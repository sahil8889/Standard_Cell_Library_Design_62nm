* File: inverter.pex.sp
* Created: Tue Dec  3 02:13:56 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt inverter  GND! OUT VDD! IN
* 
XD0_noxref GND! VDD! DIODENWX  AREA=3.6867e-12 PERIM=8.364e-06
XMMN0 OUT IN GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.3832e-13 AS=1.4144e-13
+ PD=1.572e-06 PS=1.584e-06 NRD=0.244231 NRS=0.261538 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=2.72e-07 SB=2.66e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMP0 OUT IN VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.9152e-13 AS=1.9584e-13
+ PD=1.972e-06 PS=1.984e-06 NRD=0.179167 NRS=0.188889 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=2.72e-07 SB=2.66e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=3.744e-14 PANW7=5.184e-14 PANW8=9.114e-15
+ PANW9=2.8148e-14 PANW10=4.7926e-14
*
.include "inverter.pex.sp.INVERTER.pxi"
*
.ends
*
*
