* File: AOI21.pex.sp
* Created: Mon Dec  2 22:26:54 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt AOI21  GND! OUT VDD! B A C
* 
XD0_noxref GND! VDD! DIODENWX  AREA=6.39787e-12 PERIM=1.0198e-05
XMMN2 NET18 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.5912e-13
+ PD=9.7e-07 PS=1.652e-06 NRD=0.432692 NRS=0.223077 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14
+ PANW10=0
XMMN1 OUT A NET18 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.359615 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14 PANW10=0
XMMN0 OUT C GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.5184e-13
+ PD=9.7e-07 PS=1.624e-06 NRD=0.505769 NRS=0.230769 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14
+ PANW10=0
XMMP1 NET09 B VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.2032e-13 AS=1.62e-13
+ PD=2.052e-06 PS=1.17e-06 NRD=0.141667 NRS=0.313889 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=3.744e-14 PANW7=7.2e-15 PANW8=0 PANW9=4.0362e-14
+ PANW10=9.3558e-14
XMMP0 NET09 A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.315278 NRS=0.311111 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.29642e-13 PANW10=4.8918e-14
XMMP2 OUT C NET09 VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.1024e-13 AS=1.62e-13
+ PD=2.024e-06 PS=1.17e-06 NRD=0.180556 NRS=0.309722 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=2.88e-15 PANW7=4.176e-14 PANW8=0 PANW9=4.0362e-14
+ PANW10=9.3558e-14
*
.include "AOI21.pex.sp.AOI21.pxi"
*
.ends
*
*
