* File: OAI22.pex.sp
* Created: Tue Dec  3 01:32:41 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt OAI22  GND! OUT VDD! B D C A
* 
XD0_noxref GND! VDD! DIODENWX  AREA=8.05423e-12 PERIM=1.1352e-05
XMMN0 NET12 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.5912e-13 AS=1.17e-13
+ PD=1.652e-06 PS=9.7e-07 NRD=0.192308 NRS=0.434615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14
+ PANW10=0
XMMN1 NET12 D GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.426923 NRS=0.430769 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14 PANW10=0
XMMN3 OUT C NET12 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.198077 NRS=0.438462 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14 PANW10=0
XMMN2 OUT A NET12 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.6328e-13
+ PD=9.7e-07 PS=1.668e-06 NRD=0.667308 NRS=0.223077 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14
+ PANW10=0
XMMP3 NET26 B VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2032e-13
+ PD=1.17e-06 PS=2.052e-06 NRD=0.3125 NRS=0.15 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=3.744e-14 PANW7=7.2e-15 PANW8=9.486e-15 PANW9=3.255e-14
+ PANW10=4.7244e-14
XMMP1 OUT D NET26 VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.330556 NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=9.486e-15 PANW9=7.719e-14 PANW10=9.1884e-14
XMMP0 OUT C NET27 VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.294444 NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=9.486e-15 PANW9=7.719e-14 PANW10=9.1884e-14
XMMP2 NET27 A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2608e-13
+ PD=1.17e-06 PS=2.068e-06 NRD=0.3125 NRS=0.198611 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.464e-14 PANW8=9.486e-15 PANW9=3.255e-14
+ PANW10=4.7244e-14
c_7 NET12 0 4.50891e-20
c_27 VDD! 0 4.50891e-20
*
.include "OAI22.pex.sp.OAI22.pxi"
*
.ends
*
*
