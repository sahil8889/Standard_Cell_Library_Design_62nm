* SPICE NETLIST
***************************************

.SUBCKT efuse in out
.ENDS
***************************************
.SUBCKT subc SUBCON sub
.ENDS
***************************************
.SUBCKT sblkndres IN OUT SUB
.ENDS
***************************************
.SUBCKT sblkpdres IN OUT SUB
.ENDS
***************************************
.SUBCKT esdscr_dw pd nw sx nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_tw pd nw pw nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_dw_rf pd nw sx nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_tw_rf pd nw pw nd tds1 tds2
.ENDS
***************************************
.SUBCKT npolyf_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT npolyf_u PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT ppolyf_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT nplus_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pplus_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pplus_u PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT nwella PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT indp out in gnd
.ENDS
***************************************
.SUBCKT symindp outpr outse ct BULK
.ENDS
***************************************
.SUBCKT bondpad in gp sub
.ENDS
***************************************
.SUBCKT singlecpw va vb vshield
.ENDS
***************************************
.SUBCKT coupledcpw va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT singlewire va vb vshield
.ENDS
***************************************
.SUBCKT coupledwires va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT rfline in out gnd
.ENDS
***************************************
.SUBCKT OAI22 GND! OUT VDD! B D C A
** N=39 EP=7 IP=0 FDC=9
D0 GND! VDD! diodenwx AREA=8.05423e-12 perim=1.1352e-05 $X=-26 $Y=0 $D=0
M1 GND! B 18 GND! nfet L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.5912e-13 PD=9.7e-07 PS=1.652e-06 NRD=0.434615 NRS=0.192308 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=3.06e-07 sb=1.85e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=4.774e-15 panw8=1.24e-14 panw9=1.5066e-14 panw10=0 $X=522 $Y=-1243 $D=176
M2 18 D GND! GND! nfet L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.426923 NRS=0.430769 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=8.18e-07 sb=1.338e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=4.774e-15 panw8=1.24e-14 panw9=1.5066e-14 panw10=0 $X=1034 $Y=-1243 $D=176
M3 OUT C 18 GND! nfet L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.198077 NRS=0.438462 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=1.33e-06 sb=8.26e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=4.774e-15 panw8=1.24e-14 panw9=1.5066e-14 panw10=0 $X=1546 $Y=-1243 $D=176
M4 18 A OUT GND! nfet L=6.2e-08 W=5.2e-07 AD=1.6328e-13 AS=1.17e-13 PD=1.668e-06 PS=9.7e-07 NRD=0.223077 NRS=0.667308 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=1.842e-06 sb=3.14e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=4.774e-15 panw8=1.24e-14 panw9=1.5066e-14 panw10=0 $X=2058 $Y=-1243 $D=176
M5 22 B VDD! VDD! pfet L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2032e-13 PD=1.17e-06 PS=2.052e-06 NRD=0.3125 NRS=0.15 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=3.06e-07 sb=1.85e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.744e-14 panw7=7.2e-15 panw8=9.486e-15 panw9=3.255e-14 panw10=4.7244e-14 $X=522 $Y=847 $D=189
M6 OUT D 22 VDD! pfet L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06 NRD=0.330556 NRS=0.3125 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=8.18e-07 sb=1.338e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=9.486e-15 panw9=7.719e-14 panw10=9.1884e-14 $X=1034 $Y=847 $D=189
M7 23 C OUT VDD! pfet L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06 NRD=0.3125 NRS=0.294444 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=1.33e-06 sb=8.26e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=9.486e-15 panw9=7.719e-14 panw10=9.1884e-14 $X=1546 $Y=847 $D=189
M8 VDD! A 23 VDD! pfet L=6.2e-08 W=7.2e-07 AD=2.2608e-13 AS=1.62e-13 PD=2.068e-06 PS=1.17e-06 NRD=0.198611 NRS=0.3125 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=1.842e-06 sb=3.14e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=4.464e-14 panw8=9.486e-15 panw9=3.255e-14 panw10=4.7244e-14 $X=2058 $Y=847 $D=189
.ENDS
***************************************
