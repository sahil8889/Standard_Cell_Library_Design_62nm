* SPICE NETLIST
***************************************

.SUBCKT efuse in out
.ENDS
***************************************
.SUBCKT subc SUBCON sub
.ENDS
***************************************
.SUBCKT sblkndres IN OUT SUB
.ENDS
***************************************
.SUBCKT sblkpdres IN OUT SUB
.ENDS
***************************************
.SUBCKT esdscr_dw pd nw sx nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_tw pd nw pw nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_dw_rf pd nw sx nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_tw_rf pd nw pw nd tds1 tds2
.ENDS
***************************************
.SUBCKT npolyf_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT npolyf_u PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT ppolyf_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT nplus_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pplus_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pplus_u PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT nwella PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT indp out in gnd
.ENDS
***************************************
.SUBCKT symindp outpr outse ct BULK
.ENDS
***************************************
.SUBCKT bondpad in gp sub
.ENDS
***************************************
.SUBCKT singlecpw va vb vshield
.ENDS
***************************************
.SUBCKT coupledcpw va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT singlewire va vb vshield
.ENDS
***************************************
.SUBCKT coupledwires va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT rfline in out gnd
.ENDS
***************************************
.SUBCKT inverter GND! OUT VDD! IN
** N=17 EP=4 IP=0 FDC=3
D0 GND! VDD! diodenwx AREA=3.6867e-12 perim=8.364e-06 $X=-26 $Y=0 $D=0
M1 OUT IN GND! GND! nfet L=6.2e-08 W=5.2e-07 AD=1.3832e-13 AS=1.4144e-13 PD=1.572e-06 PS=1.584e-06 NRD=0.244231 NRS=0.261538 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=2.72e-07 sb=2.66e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=5.58e-15 panw9=2.48e-14 panw10=1.86e-15 $X=522 $Y=-1430 $D=176
M2 OUT IN VDD! VDD! pfet L=6.2e-08 W=7.2e-07 AD=1.9152e-13 AS=1.9584e-13 PD=1.972e-06 PS=1.984e-06 NRD=0.179167 NRS=0.188889 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=2.72e-07 sb=2.66e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=3.744e-14 panw7=5.184e-14 panw8=9.114e-15 panw9=2.8148e-14 panw10=4.7926e-14 $X=522 $Y=853 $D=189
.ENDS
***************************************
