* File: /home/eng/s/sxv240035/cad/gf65/tutorial/AOI22/HSPICE/AOI22.pex.sp
* Created: Thu Dec  5 19:18:31 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "AOI22.pex.sp.pex"
.subckt AOI22  VSS OUT VDD B A C D
* 
* D	D
* C	C
* A	A
* B	B
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.42555e-11
+ PERIM=1.5664e-05
XMMN0 NET25 N_B_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.5756e-13 PD=9.7e-07 PS=1.646e-06 NRD=0.432692
+ NRS=0.223077 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.03e-07
+ SB=1.853e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN2 N_OUT_MMN2_d N_A_MMN2_g NET25 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.411538
+ NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=8.15e-07
+ SB=1.341e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN3 N_OUT_MMN2_d N_C_MMN3_g NET24 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.453846
+ NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.327e-06
+ SB=8.29e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN1 NET24 N_D_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.6484e-13 PD=9.7e-07 PS=1.674e-06 NRD=0.432692
+ NRS=0.225 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.839e-06
+ SB=3.17e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP3 N_NET26_MMP3_d N_B_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=2.2032e-13 AS=1.62e-13 PD=2.052e-06 PS=1.17e-06
+ NRD=0.15 NRS=0.4375 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07
+ SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
XMMP2 N_NET26_MMP2_d N_A_MMP2_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06
+ NRD=0.334722 NRS=0.1875 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15
+ PANW10=1.7608e-14
XMMP0 N_OUT_MMP0_d N_C_MMP0_g N_NET26_MMP2_d N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06 NRD=0.152778
+ NRS=0.290278 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06
+ SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.7608e-14
XMMP1 N_OUT_MMP0_d N_D_MMP1_g N_NET26_MMP1_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=2.2608e-13 PD=1.17e-06 PS=2.068e-06 NRD=0.472222
+ NRS=0.197222 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.842e-06
+ SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
*
.include "AOI22.pex.sp.AOI22.pxi"
*
.ends
*
*
