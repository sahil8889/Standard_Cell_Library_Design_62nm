* File: NAND2.pex.sp
* Created: Mon Dec  2 23:15:41 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt NAND2  GND! OUT VDD! B A
* 
XD0_noxref GND! VDD! DIODENWX  AREA=5.25006e-12 PERIM=9.414e-06
XMMN1 NET16 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.0114e-13 AS=1.5912e-13
+ PD=9.09e-07 PS=1.652e-06 NRD=0.374038 NRS=0.261538 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=7.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=1.1966e-14 PANW9=2.0274e-14 PANW10=0
XMMN0 OUT A NET16 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.43e-13 AS=1.0114e-13
+ PD=1.59e-06 PS=9.09e-07 NRD=0.217308 NRS=0.374038 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=7.57e-07 SB=2.75e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=1.1966e-14 PANW9=2.0274e-14 PANW10=0
XMMP0 OUT B VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.2032e-13 AS=1.4004e-13
+ PD=2.052e-06 PS=1.109e-06 NRD=0.188889 NRS=0.258333 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=7.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=3.744e-14 PANW7=7.2e-15 PANW8=9.114e-15 PANW9=7.4524e-14
+ PANW10=4.7926e-14
XMMP1 OUT A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.98e-13 AS=1.4004e-13
+ PD=1.99e-06 PS=1.109e-06 NRD=0.154167 NRS=0.281944 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=7.57e-07 SB=2.75e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=3.24e-14 PANW8=2.2074e-14 PANW9=7.3804e-14
+ PANW10=4.7926e-14
*
.include "NAND2.pex.sp.NAND2.pxi"
*
.ends
*
*
