* File: /home/eng/s/sxv240035/cad/gf65/tutorial/OAI21/HSPICE/OAI21.pex.sp
* Created: Thu Dec  5 19:50:51 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "OAI21.pex.sp.pex"
.subckt OAI21  VSS OUT VDD A B C
* 
* C	C
* B	B
* A	A
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.12548e-11
+ PERIM=1.3578e-05
XMMN N_NET014_MMN_d N_A_MMN_g N_VSS_MMN_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.5912e-13 AS=1.17e-13 PD=1.652e-06 PS=9.7e-07 NRD=0.192308
+ NRS=0.605769 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07
+ SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN0 N_NET014_MMN0_d N_B_MMN0_g N_VSS_MMN_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.361538
+ NRS=0.259615 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07
+ SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN1 N_OUT_MMN1_d N_C_MMN1_g N_NET014_MMN0_d N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.5184e-13 AS=1.17e-13 PD=1.624e-06 PS=9.7e-07
+ NRD=0.225 NRS=0.503846 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP1 NET19 N_A_MMP1_g N_VDD_MMP1_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=2.2032e-13 PD=1.17e-06 PS=2.052e-06 NRD=0.3125
+ NRS=0.15 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07
+ SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
XMMP0 N_OUT_MMP0_d N_B_MMP0_g NET19 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06 NRD=0.302778
+ NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07
+ SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2968e-14
XMMP2 N_OUT_MMP0_d N_C_MMP2_g N_VDD_MMP2_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=2.1024e-13 PD=1.17e-06 PS=2.024e-06 NRD=0.322222
+ NRS=0.191667 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06
+ SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=5.3902e-14 PANW10=1.8328e-14
*
.include "OAI21.pex.sp.OAI21.pxi"
*
.ends
*
*
