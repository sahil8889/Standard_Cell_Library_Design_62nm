* SPICE NETLIST
***************************************

.SUBCKT efuse in out
.ENDS
***************************************
.SUBCKT subc SUBCON sub
.ENDS
***************************************
.SUBCKT sblkndres IN OUT SUB
.ENDS
***************************************
.SUBCKT sblkpdres IN OUT SUB
.ENDS
***************************************
.SUBCKT esdscr_dw pd nw sx nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_tw pd nw pw nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_dw_rf pd nw sx nd tds1 tds2
.ENDS
***************************************
.SUBCKT esdscr_tw_rf pd nw pw nd tds1 tds2
.ENDS
***************************************
.SUBCKT npolyf_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT npolyf_u PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT ppolyf_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT nplus_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pplus_s PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT pplus_u PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT nwella PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT indp out in gnd
.ENDS
***************************************
.SUBCKT symindp outpr outse ct BULK
.ENDS
***************************************
.SUBCKT bondpad in gp sub
.ENDS
***************************************
.SUBCKT singlecpw va vb vshield
.ENDS
***************************************
.SUBCKT coupledcpw va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT singlewire va vb vshield
.ENDS
***************************************
.SUBCKT coupledwires va1 va2 vb1 vb2 vshield
.ENDS
***************************************
.SUBCKT rfline in out gnd
.ENDS
***************************************
.SUBCKT NOR3 GND! OUT VDD! A B C
** N=31 EP=6 IP=0 FDC=7
D0 GND! VDD! diodenwx AREA=6.96652e-12 perim=1.0708e-05 $X=-26 $Y=0 $D=0
M1 OUT A GND! GND! nfet L=6.2e-08 W=7e-07 AD=1.575e-13 AS=2.142e-13 PD=1.15e-06 PS=2.012e-06 NRD=0.455714 NRS=0.142857 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=3.06e-07 sb=1.316e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.2028e-14 panw10=3.1372e-14 $X=522 $Y=-1906 $D=176
M2 GND! B OUT GND! nfet L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.575e-13 PD=1.15e-06 PS=1.15e-06 NRD=0.264286 NRS=0.187143 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=8.18e-07 sb=8.04e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.2028e-14 panw10=3.1372e-14 $X=1034 $Y=-1906 $D=176
M3 OUT C GND! GND! nfet L=6.2e-08 W=7e-07 AD=2.044e-13 AS=1.575e-13 PD=1.984e-06 PS=1.15e-06 NRD=0.175714 NRS=0.378571 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=0 sa=1.33e-06 sb=2.92e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=0 panw6=0 panw7=0 panw8=0 panw9=1.2028e-14 panw10=3.1372e-14 $X=1546 $Y=-1906 $D=176
M4 17 A VDD! VDD! pfet L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=3.978e-13 PD=1.75e-06 PS=3.212e-06 NRD=0.173077 NRS=0.0830769 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=3.06e-07 sb=1.316e-06 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.1e-16 panw6=7.38e-14 panw7=2.54e-14 panw8=1.24e-14 panw9=2.9202e-14 panw10=1.4229e-13 $X=522 $Y=1329 $D=189
M5 18 B 17 VDD! pfet L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=2.925e-13 PD=1.75e-06 PS=1.75e-06 NRD=0.173077 NRS=0.173077 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=8.18e-07 sb=8.04e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.1e-16 panw6=6.2e-15 panw7=1.24e-14 panw8=1.24e-14 panw9=1.90402e-13 panw10=6.169e-14 $X=1034 $Y=1329 $D=189
M6 OUT C 18 VDD! pfet L=6.2e-08 W=1.3e-06 AD=3.796e-13 AS=2.925e-13 PD=3.184e-06 PS=1.75e-06 NRD=0.103846 NRS=0.173077 m=1 nf=1 cnr_switch=0 pccrit=0 par=1 ptwell=1 sa=1.33e-06 sb=2.92e-07 sd=0 panw1=0 panw2=0 panw3=0 panw4=0 panw5=3.1e-16 panw6=1.14e-14 panw7=8.78e-14 panw8=1.24e-14 panw9=2.9202e-14 panw10=1.4229e-13 $X=1546 $Y=1329 $D=189
.ENDS
***************************************
