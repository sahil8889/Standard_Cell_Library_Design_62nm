NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

DIVIDERCHAR "/" ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.042 ;
  SPACING 0.09 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M1

LAYER V1
  TYPE CUT ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M2

LAYER V2
  TYPE CUT ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M3

LAYER V3
  TYPE CUT ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M4

LAYER V4
  TYPE CUT ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M5

LAYER V5
  TYPE CUT ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
  END M6

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

SPACING
  SAMENET M1  M1    0.09 STACK ;
  SAMENET M2  M2    0.1 STACK ;
  SAMENET M3  M3    0.1 STACK ;
  SAMENET M4  M4    0.1 STACK ;
  SAMENET M5  M5    0.1 STACK ;
  SAMENET M6  M6    0.1 STACK ;
  SAMENET V1  V1    0.1 ;
  SAMENET V2  V2    0.1 ;
  SAMENET V3  V3    0.1 ;
  SAMENET V4  V4    0.1 ;
  SAMENET V5  V5    0.1 ;
  SAMENET V1  V2    0.00 STACK ;
  SAMENET V2  V3    0.00 STACK ;
  SAMENET V3  V4    0.00 STACK ;
  SAMENET V4  V5    0.00 STACK ;
  SAMENET V1  V3    0.00 STACK ;
  SAMENET V2  V4    0.00 STACK ;
  SAMENET V3  V5    0.00 STACK ;
  SAMENET V1  V4    0.00 STACK ;
  SAMENET V2  V5    0.00 STACK ;
  SAMENET V1  V5    0.00 STACK ;
END SPACING


VIA via5 DEFAULT
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5

VIA via4 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4

VIA via3 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3

VIA via2 DEFAULT
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2

VIA via1 DEFAULT
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1


VIARULE via1Array GENERATE
  LAYER M1 ;
  DIRECTION HORIZONTAL ;
  OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via1Array


VIARULE via2Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via2Array


VIARULE via3Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via5Array

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
  LAYER M5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
END TURNM6


SITE  CoreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 4.5 ;
END  CoreSite

SITE  TDCoverSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  TDCoverSite

SITE  SBlockSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  SBlockSite

SITE  PortCellSite
    CLASS       PAD ;
    SIZE        0.0500 BY 0.0500 ;
END  PortCellSite

SITE  Core
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 4.5 ;
END  Core

MACRO AOI21
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN AOI21 -0.026 -1.823 ;
  SIZE 2.23 BY 4.692 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.85 -0.235 0.997 0.13 ;
      LAYER M2 ;
        RECT 0.841 -0.338 0.997 0.267 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.362 -0.235 1.509 0.13 ;
      LAYER M2 ;
        RECT 1.353 -0.338 1.509 0.267 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.665 -0.503 1.817 1.76 ;
        RECT 1.207 -0.503 1.817 -0.379 ;
        RECT 1.207 -1.43 1.359 -0.379 ;
      LAYER M2 ;
        RECT 1.664 -0.338 1.82 0.267 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.08 -1.688 ;
        RECT 1.651 -1.823 1.808 -0.723 ;
        RECT 0.34 -1.823 0.497 -0.723 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.08 2.677 ;
        RECT 0.738 1.04 0.883 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.232 0.795 1.4 1.76 ;
      RECT 0.343 0.795 0.485 1.76 ;
      RECT 0.343 0.795 1.4 0.942 ;
  END
  
END AOI21

MACRO AOI22
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN AOI22 -0.026 -1.823 ;
  SIZE 2.86 BY 4.684 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.85 -0.235 0.997 0.13 ;
      LAYER M2 ;
        RECT 0.841 -0.338 0.997 0.267 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.362 -0.235 1.509 0.13 ;
      LAYER M2 ;
        RECT 1.353 -0.338 1.509 0.267 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.157 -0.235 2.304 0.13 ;
      LAYER M2 ;
        RECT 2.157 -0.338 2.313 0.267 ;
      LAYER V1 ;
        RECT 2.174 -0.05 2.274 0.05 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.635 -0.56 1.787 1.295 ;
        RECT 1.242 -0.56 1.787 -0.381 ;
        RECT 1.242 -1.379 1.394 -0.381 ;
      LAYER M2 ;
        RECT 1.63 -0.338 1.786 0.267 ;
      LAYER V1 ;
        RECT 1.641 -0.05 1.741 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.6 -1.688 ;
        RECT 2.168 -1.823 2.31 -0.723 ;
        RECT 0.343 -1.823 0.485 -0.723 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.6 2.677 ;
        RECT 0.822 0.575 0.979 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.257 2.037 2.338 2.217 ;
      RECT 2.186 0.575 2.338 2.217 ;
      RECT 1.257 0.303 1.414 2.217 ;
      RECT 0.336 0.303 0.488 1.295 ;
      RECT 0.336 0.303 1.414 0.482 ;
  END
  
END AOI22

MACRO Filler
  CLASS CORE ;
  ORIGIN 0 1.823 ;
  FOREIGN Filler 0 -1.823 ;
  SIZE 0.26 BY 4.5 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.05 -1.823 0.335 -1.688 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.05 2.549 0.335 2.677 ;
    END
  END VDD!
  
END Filler

MACRO MUX21
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN MUX21 -0.026 -1.823 ;
  SIZE 3.386 BY 4.704 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.133 -0.235 1.28 0.13 ;
      LAYER M2 ;
        RECT 1.133 -0.338 1.289 0.267 ;
      LAYER V1 ;
        RECT 1.15 -0.05 1.25 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.156 -0.235 2.303 0.13 ;
      LAYER M2 ;
        RECT 2.156 -0.338 2.312 0.267 ;
      LAYER V1 ;
        RECT 2.173 -0.05 2.273 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.681 -0.97 2.833 1.202 ;
      LAYER M2 ;
        RECT 2.681 -0.338 2.837 0.267 ;
      LAYER V1 ;
        RECT 2.696 -0.05 2.796 0.05 ;
    END
  END OUT
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.621 -0.235 0.768 0.13 ;
      LAYER M2 ;
        RECT 0.621 -0.338 0.777 0.267 ;
      LAYER V1 ;
        RECT 0.638 -0.05 0.738 0.05 ;
    END
  END S
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 3.12 -1.688 ;
        RECT 2.258 -1.823 2.4 -0.45 ;
        RECT 0.727 -1.823 0.869 -0.45 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 3.12 2.677 ;
        RECT 2.244 0.406 2.401 2.677 ;
        RECT 0.822 0.406 0.979 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.665 -1.546 1.819 1.202 ;
      RECT 0.346 -1.472 0.486 2.011 ;
  END
  
END MUX21

MACRO Merged_Cell
  CLASS CORE ;
  ORIGIN -34.32 1.823 ;
  FOREIGN Merged_Cell 34.32 -1.823 ;
  SIZE 0.26 BY 4.5 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.89 -0.235 2.037 0.13 ;
      LAYER M2 ;
        RECT 1.881 -0.338 2.037 0.267 ;
      LAYER V1 ;
        RECT 1.92 -0.05 2.02 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 17.49 -0.235 17.637 0.13 ;
      LAYER M2 ;
        RECT 17.481 -0.338 17.637 0.267 ;
      LAYER V1 ;
        RECT 17.52 -0.05 17.62 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 22.162 -0.235 22.309 0.13 ;
      LAYER M2 ;
        RECT 22.153 -0.338 22.309 0.267 ;
      LAYER V1 ;
        RECT 22.192 -0.05 22.292 0.05 ;
    END
  END C
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 31.206 -0.107 31.392 0.121 ;
      LAYER M2 ;
        RECT 31.206 -0.14 31.392 0.14 ;
      LAYER V1 ;
        RECT 31.235 -0.05 31.335 0.05 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 21.65 -0.235 21.797 0.13 ;
      LAYER M2 ;
        RECT 21.641 -0.338 21.797 0.267 ;
      LAYER V1 ;
        RECT 21.68 -0.05 21.78 0.05 ;
    END
  END D
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 24.021 -0.235 24.168 0.13 ;
      LAYER M2 ;
        RECT 24.021 -0.338 24.177 0.267 ;
      LAYER V1 ;
        RECT 24.038 -0.05 24.138 0.05 ;
    END
  END EN
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 24.533 -0.235 24.68 0.13 ;
      LAYER M2 ;
        RECT 24.533 -0.338 24.689 0.267 ;
      LAYER V1 ;
        RECT 24.55 -0.05 24.65 0.05 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 27.89 -0.512 28.058 1.308 ;
        RECT 27.481 -0.512 28.058 -0.388 ;
        RECT 27.481 -1.127 27.633 -0.388 ;
      LAYER M2 ;
        RECT 27.89 -0.338 28.058 0.267 ;
      LAYER V1 ;
        RECT 27.925 -0.05 28.025 0.05 ;
    END
  END OUT
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 32.098 -0.952 32.215 1.157 ;
      LAYER M2 ;
        RECT 32.029 -0.14 32.215 0.14 ;
      LAYER V1 ;
        RECT 32.104 -0.05 32.204 0.05 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 30.147 -0.107 30.333 0.121 ;
      LAYER M2 ;
        RECT 30.147 -0.14 30.333 0.14 ;
      LAYER V1 ;
        RECT 30.194 -0.05 30.294 0.05 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.341 -0.235 6.488 0.13 ;
      LAYER M2 ;
        RECT 6.341 -0.338 6.497 0.267 ;
      LAYER V1 ;
        RECT 6.358 -0.05 6.458 0.05 ;
    END
  END S
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 34.655 -1.688 ;
        RECT 34.074 -1.83 34.184 -0.411 ;
        RECT 33.488 -1.83 33.598 -0.411 ;
        RECT 32.521 -1.83 32.631 -0.411 ;
        RECT 31.48 -1.83 31.59 -0.411 ;
        RECT 30.729 -1.83 30.819 -0.305 ;
        RECT 30.204 -1.83 30.294 -0.328 ;
        RECT 29.188 -1.83 29.298 -0.411 ;
        RECT 28.389 -1.823 28.546 -0.607 ;
        RECT 27.078 -1.823 27.235 -0.607 ;
        RECT 26.048 -1.823 26.19 -0.607 ;
        RECT 24.127 -1.823 24.269 -0.479 ;
        RECT 21.538 -1.823 21.68 -0.723 ;
        RECT 19.542 -1.823 19.699 -0.91 ;
        RECT 17.847 -1.823 17.999 -0.91 ;
        RECT 16.983 -1.823 17.125 -0.91 ;
        RECT 15.775 -1.823 15.927 -0.91 ;
        RECT 12.823 -1.823 12.965 -0.91 ;
        RECT 10.743 -1.823 10.885 -0.91 ;
        RECT 9.148 -1.823 9.29 -0.694 ;
        RECT 7.978 -1.823 8.12 -0.45 ;
        RECT 6.447 -1.823 6.589 -0.45 ;
        RECT 5.288 -1.823 5.43 -0.723 ;
        RECT 3.463 -1.823 3.605 -0.723 ;
        RECT 2.691 -1.823 2.848 -0.723 ;
        RECT 1.38 -1.823 1.537 -0.723 ;
        RECT 0.308 -1.823 0.45 -0.73 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.001 2.549 34.655 2.677 ;
        RECT 33.493 0.41 33.593 2.677 ;
        RECT 32.527 0.41 32.627 2.677 ;
        RECT 31.32 0.41 31.42 2.677 ;
        RECT 30.155 0.441 30.255 2.677 ;
        RECT 29.194 0.441 29.294 2.677 ;
        RECT 26.959 0.588 27.101 2.677 ;
        RECT 24.222 0.351 24.379 2.677 ;
        RECT 22.986 0.847 23.138 2.677 ;
        RECT 21.136 0.524 21.288 2.677 ;
        RECT 20.388 0.853 20.54 2.677 ;
        RECT 19.063 0.853 19.208 2.677 ;
        RECT 16.976 0.853 17.128 2.677 ;
        RECT 15.39 0.853 15.547 2.677 ;
        RECT 14.666 0.853 14.818 2.677 ;
        RECT 13.814 0.853 13.971 2.677 ;
        RECT 12.816 0.853 12.968 2.677 ;
        RECT 11.607 0.853 11.759 2.677 ;
        RECT 10.736 0.853 10.888 2.677 ;
        RECT 9.535 0.853 9.687 2.677 ;
        RECT 7.964 0.406 8.121 2.677 ;
        RECT 6.542 0.406 6.699 2.677 ;
        RECT 3.942 0.575 4.099 2.677 ;
        RECT 1.778 1.04 1.923 2.677 ;
        RECT 0.31 0.853 0.467 2.677 ;
    END
  END VDD!
  PIN A_mj1
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 26.529 -0.235 26.676 0.13 ;
      LAYER M2 ;
        RECT 26.52 -0.338 26.676 0.267 ;
      LAYER V1 ;
        RECT 26.559 -0.05 26.659 0.05 ;
    END
  END A_mj1
  PIN A_mj2
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 22.957 -0.235 23.104 0.13 ;
      LAYER M2 ;
        RECT 22.957 -0.338 23.113 0.267 ;
      LAYER V1 ;
        RECT 22.974 -0.05 23.074 0.05 ;
    END
  END A_mj2
  PIN A_mj3
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 19.058 -0.235 19.205 0.13 ;
      LAYER M2 ;
        RECT 19.049 -0.338 19.205 0.267 ;
      LAYER V1 ;
        RECT 19.088 -0.05 19.188 0.05 ;
    END
  END A_mj3
  PIN A_mj4
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.978 -0.235 17.125 0.13 ;
      LAYER M2 ;
        RECT 16.969 -0.338 17.125 0.267 ;
      LAYER V1 ;
        RECT 17.008 -0.05 17.108 0.05 ;
    END
  END A_mj4
  PIN A_mj5
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 15.418 -0.235 15.565 0.13 ;
      LAYER M2 ;
        RECT 15.409 -0.338 15.565 0.267 ;
      LAYER V1 ;
        RECT 15.448 -0.05 15.548 0.05 ;
    END
  END A_mj5
  PIN A_mj6
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.354 -0.235 14.501 0.13 ;
      LAYER M2 ;
        RECT 14.345 -0.338 14.501 0.267 ;
      LAYER V1 ;
        RECT 14.384 -0.05 14.484 0.05 ;
    END
  END A_mj6
  PIN A_mj7
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.762 -0.235 11.909 0.13 ;
      LAYER M2 ;
        RECT 11.753 -0.338 11.909 0.267 ;
      LAYER V1 ;
        RECT 11.792 -0.05 11.892 0.05 ;
    END
  END A_mj7
  PIN A_mj8
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.629 -0.235 9.776 0.13 ;
      LAYER M2 ;
        RECT 9.62 -0.338 9.776 0.267 ;
      LAYER V1 ;
        RECT 9.659 -0.05 9.759 0.05 ;
    END
  END A_mj8
  PIN A_mj9
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.853 -0.235 7 0.13 ;
      LAYER M2 ;
        RECT 6.853 -0.338 7.009 0.267 ;
      LAYER V1 ;
        RECT 6.87 -0.05 6.97 0.05 ;
    END
  END A_mj9
  PIN A_mj10
    MUSTJOIN A ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.97 -0.235 4.117 0.13 ;
      LAYER M2 ;
        RECT 3.961 -0.338 4.117 0.267 ;
      LAYER V1 ;
        RECT 4 -0.05 4.1 0.05 ;
    END
  END A_mj10
  PIN B_mj1
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.378 -0.235 1.525 0.13 ;
      LAYER M2 ;
        RECT 1.369 -0.338 1.525 0.267 ;
      LAYER V1 ;
        RECT 1.408 -0.05 1.508 0.05 ;
    END
  END B_mj1
  PIN B_mj2
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.458 -0.235 3.605 0.13 ;
      LAYER M2 ;
        RECT 3.449 -0.338 3.605 0.267 ;
      LAYER V1 ;
        RECT 3.488 -0.05 3.588 0.05 ;
    END
  END B_mj2
  PIN B_mj3
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.876 -0.235 8.023 0.13 ;
      LAYER M2 ;
        RECT 7.876 -0.338 8.032 0.267 ;
      LAYER V1 ;
        RECT 7.893 -0.05 7.993 0.05 ;
    END
  END B_mj3
  PIN B_mj4
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.178 -0.235 9.325 0.13 ;
      LAYER M2 ;
        RECT 9.169 -0.338 9.325 0.267 ;
      LAYER V1 ;
        RECT 9.208 -0.05 9.308 0.05 ;
    END
  END B_mj4
  PIN B_mj5
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.25 -0.235 11.397 0.13 ;
      LAYER M2 ;
        RECT 11.241 -0.338 11.397 0.267 ;
      LAYER V1 ;
        RECT 11.28 -0.05 11.38 0.05 ;
    END
  END B_mj5
  PIN B_mj6
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.842 -0.235 13.989 0.13 ;
      LAYER M2 ;
        RECT 13.833 -0.338 13.989 0.267 ;
      LAYER V1 ;
        RECT 13.872 -0.05 13.972 0.05 ;
    END
  END B_mj6
  PIN B_mj7
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 15.869 -0.235 16.016 0.13 ;
      LAYER M2 ;
        RECT 15.86 -0.338 16.016 0.267 ;
      LAYER V1 ;
        RECT 15.899 -0.05 15.999 0.05 ;
    END
  END B_mj7
  PIN B_mj8
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 19.57 -0.235 19.717 0.13 ;
      LAYER M2 ;
        RECT 19.561 -0.338 19.717 0.267 ;
      LAYER V1 ;
        RECT 19.6 -0.05 19.7 0.05 ;
    END
  END B_mj8
  PIN B_mj9
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 21.138 -0.235 21.285 0.13 ;
      LAYER M2 ;
        RECT 21.129 -0.338 21.285 0.267 ;
      LAYER V1 ;
        RECT 21.168 -0.05 21.268 0.05 ;
    END
  END B_mj9
  PIN B_mj10
    MUSTJOIN B ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 26.078 -0.235 26.225 0.13 ;
      LAYER M2 ;
        RECT 26.069 -0.338 26.225 0.267 ;
      LAYER V1 ;
        RECT 26.108 -0.05 26.208 0.05 ;
    END
  END B_mj10
  PIN C_mj1
    MUSTJOIN C ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 20.082 -0.235 20.229 0.13 ;
      LAYER M2 ;
        RECT 20.073 -0.338 20.229 0.267 ;
      LAYER V1 ;
        RECT 20.112 -0.05 20.212 0.05 ;
    END
  END C_mj1
  PIN C_mj2
    MUSTJOIN C ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.402 -0.235 2.549 0.13 ;
      LAYER M2 ;
        RECT 2.393 -0.338 2.549 0.267 ;
      LAYER V1 ;
        RECT 2.432 -0.05 2.532 0.05 ;
    END
  END C_mj2
  PIN C_mj3
    MUSTJOIN C ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 18.002 -0.235 18.149 0.13 ;
      LAYER M2 ;
        RECT 17.993 -0.338 18.149 0.267 ;
      LAYER V1 ;
        RECT 18.032 -0.05 18.132 0.05 ;
    END
  END C_mj3
  PIN C_mj4
    MUSTJOIN C ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.33 -0.235 13.477 0.13 ;
      LAYER M2 ;
        RECT 13.321 -0.338 13.477 0.267 ;
      LAYER V1 ;
        RECT 13.36 -0.05 13.46 0.05 ;
    END
  END C_mj4
  PIN C_mj5
    MUSTJOIN C ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.482 -0.235 4.629 0.13 ;
      LAYER M2 ;
        RECT 4.473 -0.338 4.629 0.267 ;
      LAYER V1 ;
        RECT 4.512 -0.05 4.612 0.05 ;
    END
  END C_mj5
  PIN C_mj6
    MUSTJOIN C ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.738 -0.235 10.885 0.13 ;
      LAYER M2 ;
        RECT 10.729 -0.338 10.885 0.267 ;
      LAYER V1 ;
        RECT 10.768 -0.05 10.868 0.05 ;
    END
  END C_mj6
  PIN D_mj1
    MUSTJOIN D ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 29.141 -0.107 29.327 0.121 ;
      LAYER M2 ;
        RECT 29.141 -0.14 29.327 0.14 ;
      LAYER V1 ;
        RECT 29.188 -0.05 29.288 0.05 ;
    END
  END D_mj1
  PIN D_mj2
    MUSTJOIN D ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.277 -0.235 5.424 0.13 ;
      LAYER M2 ;
        RECT 5.277 -0.338 5.433 0.267 ;
      LAYER V1 ;
        RECT 5.294 -0.05 5.394 0.05 ;
    END
  END D_mj2
  PIN D_mj3
    MUSTJOIN D ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.818 -0.235 12.965 0.13 ;
      LAYER M2 ;
        RECT 12.809 -0.338 12.965 0.267 ;
      LAYER V1 ;
        RECT 12.848 -0.05 12.948 0.05 ;
    END
  END D_mj3
  PIN IN_mj1
    MUSTJOIN IN ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END IN_mj1
  PIN OUT_mj1
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 22.057 0.529 22.586 0.708 ;
        RECT 22.434 -1.243 22.586 0.708 ;
        RECT 22.057 0.529 22.214 1.567 ;
      LAYER M2 ;
        RECT 22.43 -0.338 22.586 0.267 ;
      LAYER V1 ;
        RECT 22.441 -0.05 22.541 0.05 ;
    END
  END OUT_mj1
  PIN OUT_mj2
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 25.065 -0.999 25.217 1.071 ;
      LAYER M2 ;
        RECT 25.064 -0.338 25.22 0.267 ;
      LAYER V1 ;
        RECT 25.075 -0.05 25.175 0.05 ;
    END
  END OUT_mj2
  PIN OUT_mj3
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 19.952 0.508 20.537 0.634 ;
        RECT 20.385 -1.43 20.537 0.634 ;
        RECT 19.952 0.508 20.12 1.573 ;
      LAYER M2 ;
        RECT 20.384 -0.338 20.54 0.267 ;
      LAYER V1 ;
        RECT 20.395 -0.05 20.495 0.05 ;
    END
  END OUT_mj3
  PIN OUT_mj4
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 18.305 -1.43 18.457 1.573 ;
        RECT 17.462 -0.505 18.457 -0.379 ;
        RECT 17.462 -1.427 17.619 -0.379 ;
      LAYER M2 ;
        RECT 18.304 -0.338 18.46 0.267 ;
      LAYER V1 ;
        RECT 18.315 -0.05 18.415 0.05 ;
    END
  END OUT_mj4
  PIN OUT_mj5
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.154 -1.43 16.306 1.573 ;
        RECT 15.388 -0.577 16.306 -0.451 ;
        RECT 15.388 -1.43 15.53 -0.451 ;
      LAYER M2 ;
        RECT 16.154 -0.338 16.31 0.267 ;
      LAYER V1 ;
        RECT 16.182 -0.05 16.282 0.05 ;
    END
  END OUT_mj5
  PIN OUT_mj6
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.302 0.483 14.809 0.662 ;
        RECT 14.657 -1.43 14.809 0.662 ;
        RECT 14.199 0.483 14.351 1.573 ;
        RECT 13.302 0.483 13.459 1.573 ;
      LAYER M2 ;
        RECT 14.656 -0.338 14.812 0.267 ;
      LAYER V1 ;
        RECT 14.667 -0.05 14.767 0.05 ;
    END
  END OUT_mj6
  PIN OUT_mj7
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.065 -1.43 12.217 1.573 ;
        RECT 11.222 0.458 12.217 0.584 ;
        RECT 11.222 0.458 11.379 1.573 ;
      LAYER M2 ;
        RECT 12.064 -0.338 12.22 0.267 ;
      LAYER V1 ;
        RECT 12.075 -0.05 12.175 0.05 ;
    END
  END OUT_mj7
  PIN OUT_mj8
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.914 -1.514 10.066 1.573 ;
        RECT 9.15 0.458 10.066 0.584 ;
        RECT 9.15 0.458 9.307 1.573 ;
      LAYER M2 ;
        RECT 9.914 -0.338 10.07 0.267 ;
      LAYER V1 ;
        RECT 9.942 -0.05 10.042 0.05 ;
    END
  END OUT_mj8
  PIN OUT_mj9
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.401 -0.97 8.553 1.202 ;
      LAYER M2 ;
        RECT 8.401 -0.338 8.557 0.267 ;
      LAYER V1 ;
        RECT 8.416 -0.05 8.516 0.05 ;
    END
  END OUT_mj9
  PIN OUT_mj10
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.755 -0.56 4.907 1.295 ;
        RECT 4.362 -0.56 4.907 -0.381 ;
        RECT 4.362 -1.379 4.514 -0.381 ;
      LAYER M2 ;
        RECT 4.75 -0.338 4.906 0.267 ;
      LAYER V1 ;
        RECT 4.761 -0.05 4.861 0.05 ;
    END
  END OUT_mj10
  PIN OUT_mj11
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.705 -0.503 2.857 1.76 ;
        RECT 2.247 -0.503 2.857 -0.379 ;
        RECT 2.247 -1.43 2.399 -0.379 ;
      LAYER M2 ;
        RECT 2.704 -0.338 2.86 0.267 ;
      LAYER V1 ;
        RECT 2.715 -0.05 2.815 0.05 ;
    END
  END OUT_mj11
  PIN OUT_mj12
    MUSTJOIN OUT ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.638 -1.43 0.79 2.153 ;
      LAYER M2 ;
        RECT 0.638 -0.355 0.741 0.264 ;
      LAYER V1 ;
        RECT 0.641 -0.05 0.741 0.05 ;
    END
  END OUT_mj12
  OBS
    LAYER M1 ;
      RECT 34.075 -0.321 34.185 1.13 ;
      RECT 33.384 0.177 34.185 0.317 ;
      RECT 33.813 -0.321 34.185 -0.231 ;
      RECT 33.813 -0.931 33.923 -0.231 ;
      RECT 32.976 -0.983 33.086 1.227 ;
      RECT 32.416 0.177 33.086 0.317 ;
      RECT 32.976 -0.141 33.968 -0.001 ;
      RECT 31.741 1.256 32.187 1.346 ;
      RECT 31.741 -1.594 31.832 1.346 ;
      RECT 31.741 -1.545 32.429 -1.455 ;
      RECT 30.98 0.23 31.07 2.26 ;
      RECT 30.345 2.135 31.23 2.225 ;
      RECT 30.97 0.23 31.625 0.32 ;
      RECT 31.485 -0.321 31.625 0.32 ;
      RECT 30.971 -0.321 31.625 -0.231 ;
      RECT 30.98 -1.037 31.07 -0.231 ;
      RECT 30.729 0.031 30.819 1.561 ;
      RECT 30.051 0.211 30.829 0.351 ;
      RECT 30.456 0.031 30.829 0.121 ;
      RECT 30.456 -0.931 30.566 0.121 ;
      RECT 29.652 -1.315 29.742 1.202 ;
      RECT 29.652 -1.315 30.114 -1.225 ;
      RECT 27.476 1.954 28.555 2.101 ;
      RECT 28.403 0.588 28.555 2.101 ;
      RECT 27.476 0.588 27.621 2.101 ;
      RECT 26.05 0.363 26.207 1.308 ;
      RECT 26.05 0.363 27.223 0.489 ;
      RECT 27.076 -0.511 27.223 0.489 ;
      RECT 26.435 -0.511 27.223 -0.385 ;
      RECT 26.435 -1.303 26.587 -0.385 ;
      RECT 24.607 1.745 25.522 1.873 ;
      RECT 25.39 -1.494 25.522 1.873 ;
      RECT 24.607 0.351 24.759 1.873 ;
      RECT 24.607 -1.494 24.759 -0.479 ;
      RECT 24.607 -1.494 25.522 -1.369 ;
      RECT 21.142 -0.624 22.194 -0.478 ;
      RECT 22.042 -1.547 22.194 -0.478 ;
      RECT 21.144 -1.243 21.296 -0.478 ;
      RECT 22.968 -1.547 23.11 -0.723 ;
      RECT 22.042 -1.547 23.11 -1.401 ;
      RECT 19.063 -0.505 20.079 -0.379 ;
      RECT 19.927 -1.43 20.079 -0.379 ;
      RECT 19.063 -1.43 19.205 -0.379 ;
      RECT 4.377 2.037 5.458 2.217 ;
      RECT 5.306 0.575 5.458 2.217 ;
      RECT 4.377 0.303 4.534 2.217 ;
      RECT 3.456 0.303 3.608 1.295 ;
      RECT 3.456 0.303 4.534 0.482 ;
      RECT 2.272 0.795 2.44 1.76 ;
      RECT 1.383 0.795 1.525 1.76 ;
      RECT 1.383 0.795 2.44 0.942 ;
      RECT 32.717 2.367 33.394 2.457 ;
      RECT 31.51 1.436 32.437 1.526 ;
      RECT 31.51 1.902 32.437 1.992 ;
      RECT 31.51 2.135 32.437 2.225 ;
      RECT 31.76 2.368 32.437 2.458 ;
      RECT 31.51 1.669 31.983 1.759 ;
      RECT 30.909 -1.545 31.39 -1.455 ;
      RECT 30.35 1.669 30.89 1.759 ;
      RECT 30.345 1.902 30.831 1.992 ;
      RECT 29.597 -1.545 30.114 -1.455 ;
      RECT 23.642 -0.999 23.794 2.032 ;
      RECT 7.385 -1.546 7.539 1.202 ;
      RECT 6.066 -1.472 6.206 2.011 ;
  END
  
END Merged_Cell

MACRO NAND2
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN NAND2 -0.026 -1.823 ;
  SIZE 1.816 BY 4.714 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.789 -0.235 0.936 0.13 ;
      LAYER M2 ;
        RECT 0.78 -0.338 0.936 0.267 ;
      LAYER V1 ;
        RECT 0.819 -0.05 0.919 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.074 -1.514 1.226 1.573 ;
        RECT 0.31 0.458 1.226 0.584 ;
        RECT 0.31 0.458 0.467 1.573 ;
      LAYER M2 ;
        RECT 1.074 -0.338 1.23 0.267 ;
      LAYER V1 ;
        RECT 1.102 -0.05 1.202 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 1.56 -1.688 ;
        RECT 0.308 -1.823 0.45 -0.694 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 1.56 2.677 ;
        RECT 0.695 0.853 0.847 2.677 ;
    END
  END VDD!
  
END NAND2

MACRO NAND3
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN NAND3 -0.026 -1.823 ;
  SIZE 2.394 BY 4.671 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.362 -0.235 1.509 0.13 ;
      LAYER M2 ;
        RECT 1.353 -0.338 1.509 0.267 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.85 -0.235 0.997 0.13 ;
      LAYER M2 ;
        RECT 0.841 -0.338 0.997 0.267 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.665 -1.43 1.817 1.573 ;
        RECT 0.822 0.458 1.817 0.584 ;
        RECT 0.822 0.458 0.979 1.573 ;
      LAYER M2 ;
        RECT 1.664 -0.338 1.82 0.267 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.08 -1.688 ;
        RECT 0.343 -1.823 0.485 -0.91 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.007 2.549 2.073 2.677 ;
        RECT 1.207 0.853 1.359 2.677 ;
        RECT 0.336 0.853 0.488 2.677 ;
    END
  END VDD!
  
END NAND3

MACRO NAND4
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN NAND4 -0.026 -1.823 ;
  SIZE 2.844 BY 4.656 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.874 -0.235 2.021 0.13 ;
      LAYER M2 ;
        RECT 1.865 -0.338 2.021 0.267 ;
      LAYER V1 ;
        RECT 1.904 -0.05 2.004 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.362 -0.235 1.509 0.13 ;
      LAYER M2 ;
        RECT 1.353 -0.338 1.509 0.267 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.85 -0.235 0.997 0.13 ;
      LAYER M2 ;
        RECT 0.841 -0.338 0.997 0.267 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.822 0.483 2.329 0.662 ;
        RECT 2.177 -1.43 2.329 0.662 ;
        RECT 1.719 0.483 1.871 1.573 ;
        RECT 0.822 0.483 0.979 1.573 ;
      LAYER M2 ;
        RECT 2.176 -0.338 2.332 0.267 ;
      LAYER V1 ;
        RECT 2.187 -0.05 2.287 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.6 -1.688 ;
        RECT 0.343 -1.823 0.485 -0.91 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.6 2.677 ;
        RECT 2.186 0.853 2.338 2.677 ;
        RECT 1.334 0.853 1.491 2.677 ;
        RECT 0.336 0.853 0.488 2.677 ;
    END
  END VDD!
  
END NAND4

MACRO NOR2
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN NOR2 -0.026 -1.823 ;
  SIZE 1.832 BY 4.741 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.789 -0.235 0.936 0.13 ;
      LAYER M2 ;
        RECT 0.78 -0.338 0.936 0.267 ;
      LAYER V1 ;
        RECT 0.819 -0.05 0.919 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.074 -1.43 1.226 1.573 ;
        RECT 0.308 -0.577 1.226 -0.451 ;
        RECT 0.308 -1.43 0.45 -0.451 ;
      LAYER M2 ;
        RECT 1.074 -0.338 1.23 0.267 ;
      LAYER V1 ;
        RECT 1.102 -0.05 1.202 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 1.56 -1.688 ;
        RECT 0.695 -1.823 0.847 -0.91 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 1.56 2.677 ;
        RECT 0.31 0.853 0.467 2.677 ;
    END
  END VDD!
  
END NOR2

MACRO NOR3
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN NOR3 -0.026 -1.823 ;
  SIZE 2.369 BY 4.674 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.85 -0.235 0.997 0.13 ;
      LAYER M2 ;
        RECT 0.841 -0.338 0.997 0.267 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.362 -0.235 1.509 0.13 ;
      LAYER M2 ;
        RECT 1.353 -0.338 1.509 0.267 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.665 -1.43 1.817 1.573 ;
        RECT 0.822 -0.505 1.817 -0.379 ;
        RECT 0.822 -1.427 0.979 -0.379 ;
      LAYER M2 ;
        RECT 1.664 -0.338 1.82 0.267 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.08 -1.688 ;
        RECT 1.207 -1.823 1.359 -0.91 ;
        RECT 0.343 -1.823 0.485 -0.91 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.08 2.677 ;
        RECT 0.336 0.853 0.488 2.677 ;
    END
  END VDD!
  
END NOR3

MACRO OAI21
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN OAI21 -0.026 -1.823 ;
  SIZE 2.325 BY 4.745 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.85 -0.235 0.997 0.13 ;
      LAYER M2 ;
        RECT 0.841 -0.338 0.997 0.267 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.362 -0.235 1.509 0.13 ;
      LAYER M2 ;
        RECT 1.353 -0.338 1.509 0.267 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.232 0.508 1.817 0.634 ;
        RECT 1.665 -1.43 1.817 0.634 ;
        RECT 1.232 0.508 1.4 1.573 ;
      LAYER M2 ;
        RECT 1.664 -0.338 1.82 0.267 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.08 -1.688 ;
        RECT 0.822 -1.823 0.979 -0.91 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.08 2.677 ;
        RECT 1.668 0.853 1.82 2.677 ;
        RECT 0.343 0.853 0.488 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 0.343 -0.505 1.359 -0.379 ;
      RECT 1.207 -1.43 1.359 -0.379 ;
      RECT 0.343 -1.43 0.485 -0.379 ;
  END
  
END OAI21

MACRO OAI22
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN OAI22 -0.026 -1.823 ;
  SIZE 2.834 BY 4.665 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.157 -0.235 2.304 0.13 ;
      LAYER M2 ;
        RECT 2.157 -0.338 2.313 0.267 ;
      LAYER V1 ;
        RECT 2.174 -0.05 2.274 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.362 -0.235 1.509 0.13 ;
      LAYER M2 ;
        RECT 1.353 -0.338 1.509 0.267 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.85 -0.235 0.997 0.13 ;
      LAYER M2 ;
        RECT 0.841 -0.338 0.997 0.267 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.257 0.529 1.786 0.708 ;
        RECT 1.634 -1.243 1.786 0.708 ;
        RECT 1.257 0.529 1.414 1.567 ;
      LAYER M2 ;
        RECT 1.63 -0.338 1.786 0.267 ;
      LAYER V1 ;
        RECT 1.641 -0.05 1.741 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.6 -1.688 ;
        RECT 0.738 -1.823 0.88 -0.723 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.6 2.677 ;
        RECT 2.186 0.847 2.338 2.677 ;
        RECT 0.336 0.524 0.488 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 0.342 -0.624 1.394 -0.478 ;
      RECT 1.242 -1.547 1.394 -0.478 ;
      RECT 0.344 -1.243 0.496 -0.478 ;
      RECT 2.168 -1.547 2.31 -0.723 ;
      RECT 1.242 -1.547 2.31 -1.401 ;
  END
  
END OAI22

MACRO Tri_INV
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN Tri_INV -0.026 -1.823 ;
  SIZE 2.575 BY 4.719 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.621 -0.235 0.768 0.13 ;
      LAYER M2 ;
        RECT 0.621 -0.338 0.777 0.267 ;
      LAYER V1 ;
        RECT 0.638 -0.05 0.738 0.05 ;
    END
  END EN
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.133 -0.235 1.28 0.13 ;
      LAYER M2 ;
        RECT 1.133 -0.338 1.289 0.267 ;
      LAYER V1 ;
        RECT 1.15 -0.05 1.25 0.05 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.665 -0.999 1.817 1.071 ;
      LAYER M2 ;
        RECT 1.664 -0.338 1.82 0.267 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 2.34 -1.688 ;
        RECT 0.727 -1.823 0.869 -0.479 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.34 2.677 ;
        RECT 0.822 0.351 0.979 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.207 1.745 2.122 1.873 ;
      RECT 1.99 -1.494 2.122 1.873 ;
      RECT 1.207 0.351 1.359 1.873 ;
      RECT 1.207 -1.494 1.359 -0.479 ;
      RECT 1.207 -1.494 2.122 -1.369 ;
      RECT 0.242 -0.999 0.394 2.032 ;
  END
  
END Tri_INV

MACRO XOR2
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN XOR2 -0.026 -1.823 ;
  SIZE 3.354 BY 4.784 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.789 -0.235 0.936 0.13 ;
      LAYER M2 ;
        RECT 0.78 -0.338 0.936 0.267 ;
      LAYER V1 ;
        RECT 0.819 -0.05 0.919 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.15 -0.512 2.318 1.308 ;
        RECT 1.741 -0.512 2.318 -0.388 ;
        RECT 1.741 -1.127 1.893 -0.388 ;
      LAYER M2 ;
        RECT 2.15 -0.338 2.318 0.267 ;
      LAYER V1 ;
        RECT 2.185 -0.05 2.285 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 3.12 -1.688 ;
        RECT 2.649 -1.823 2.806 -0.607 ;
        RECT 1.338 -1.823 1.495 -0.607 ;
        RECT 0.308 -1.823 0.45 -0.607 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 3.12 2.677 ;
        RECT 1.219 0.588 1.361 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.736 1.954 2.815 2.101 ;
      RECT 2.663 0.588 2.815 2.101 ;
      RECT 1.736 0.588 1.881 2.101 ;
      RECT 0.31 0.363 0.467 1.308 ;
      RECT 0.31 0.363 1.483 0.489 ;
      RECT 1.336 -0.511 1.483 0.489 ;
      RECT 0.695 -0.511 1.483 -0.385 ;
      RECT 0.695 -1.303 0.847 -0.385 ;
  END
  
END XOR2

MACRO dff
  CLASS CORE ;
  ORIGIN 0.136 1.83 ;
  FOREIGN dff -0.136 -1.83 ;
  SIZE 5.745 BY 4.699 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.346 -0.107 2.532 0.121 ;
      LAYER M2 ;
        RECT 2.346 -0.14 2.532 0.14 ;
      LAYER V1 ;
        RECT 2.375 -0.05 2.475 0.05 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.281 -0.107 0.467 0.121 ;
      LAYER M2 ;
        RECT 0.281 -0.14 0.467 0.14 ;
      LAYER V1 ;
        RECT 0.328 -0.05 0.428 0.05 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.238 -0.952 3.355 1.157 ;
      LAYER M2 ;
        RECT 3.169 -0.14 3.355 0.14 ;
      LAYER V1 ;
        RECT 3.244 -0.05 3.344 0.05 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.287 -0.107 1.473 0.121 ;
      LAYER M2 ;
        RECT 1.287 -0.14 1.473 0.14 ;
      LAYER V1 ;
        RECT 1.334 -0.05 1.434 0.05 ;
    END
  END R
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 5.46 -1.688 ;
        RECT 5.214 -1.83 5.324 -0.411 ;
        RECT 4.628 -1.83 4.738 -0.411 ;
        RECT 3.661 -1.83 3.771 -0.411 ;
        RECT 2.62 -1.83 2.73 -0.411 ;
        RECT 1.869 -1.83 1.959 -0.305 ;
        RECT 1.344 -1.83 1.434 -0.328 ;
        RECT 0.328 -1.83 0.438 -0.411 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 5.46 2.677 ;
        RECT 4.633 0.41 4.733 2.677 ;
        RECT 3.667 0.41 3.767 2.677 ;
        RECT 2.46 0.41 2.56 2.677 ;
        RECT 1.295 0.441 1.395 2.677 ;
        RECT 0.334 0.441 0.434 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 5.215 -0.321 5.325 1.13 ;
      RECT 4.524 0.177 5.325 0.317 ;
      RECT 4.953 -0.321 5.325 -0.231 ;
      RECT 4.953 -0.931 5.063 -0.231 ;
      RECT 4.116 -0.983 4.226 1.227 ;
      RECT 3.556 0.177 4.226 0.317 ;
      RECT 4.116 -0.141 5.108 -0.001 ;
      RECT 2.881 1.256 3.327 1.346 ;
      RECT 2.881 -1.594 2.972 1.346 ;
      RECT 2.881 -1.545 3.569 -1.455 ;
      RECT 2.12 0.23 2.21 2.26 ;
      RECT 1.485 2.135 2.37 2.225 ;
      RECT 2.11 0.23 2.765 0.32 ;
      RECT 2.625 -0.321 2.765 0.32 ;
      RECT 2.111 -0.321 2.765 -0.231 ;
      RECT 2.12 -1.037 2.21 -0.231 ;
      RECT 1.869 0.031 1.959 1.561 ;
      RECT 1.191 0.211 1.969 0.351 ;
      RECT 1.596 0.031 1.969 0.121 ;
      RECT 1.596 -0.931 1.706 0.121 ;
      RECT 0.792 -1.315 0.882 1.202 ;
      RECT 0.792 -1.315 1.254 -1.225 ;
      RECT 3.857 2.367 4.534 2.457 ;
      RECT 2.65 1.436 3.577 1.526 ;
      RECT 2.65 1.902 3.577 1.992 ;
      RECT 2.65 2.135 3.577 2.225 ;
      RECT 2.9 2.368 3.577 2.458 ;
      RECT 2.65 1.669 3.123 1.759 ;
      RECT 2.049 -1.545 2.53 -1.455 ;
      RECT 1.49 1.669 2.03 1.759 ;
      RECT 1.485 1.902 1.971 1.992 ;
      RECT 0.737 -1.545 1.254 -1.455 ;
  END
  
END dff

MACRO inverter
  CLASS CORE ;
  ORIGIN 0.026 1.823 ;
  FOREIGN inverter -0.026 -1.823 ;
  SIZE 1.263 BY 4.742 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.338 -0.235 0.485 0.13 ;
      LAYER M2 ;
        RECT 0.329 -0.338 0.485 0.267 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.638 -1.43 0.79 2.153 ;
      LAYER M2 ;
        RECT 0.638 -0.355 0.741 0.264 ;
      LAYER V1 ;
        RECT 0.641 -0.05 0.741 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 1.04 -1.688 ;
        RECT 0.308 -1.823 0.45 -0.73 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.001 2.549 1.04 2.677 ;
        RECT 0.31 0.853 0.467 2.677 ;
    END
  END VDD!
  
END inverter

END LIBRARY
