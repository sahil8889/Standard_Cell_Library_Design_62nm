NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

DIVIDERCHAR "/" ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.042 ;
  SPACING 0.09 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M1

LAYER V1
  TYPE CUT ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M2

LAYER V2
  TYPE CUT ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M3

LAYER V3
  TYPE CUT ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M4

LAYER V4
  TYPE CUT ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M5

LAYER V5
  TYPE CUT ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
  END M6

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

SPACING
  SAMENET M1  M1    0.09 STACK ;
  SAMENET M2  M2    0.1 STACK ;
  SAMENET M3  M3    0.1 STACK ;
  SAMENET M4  M4    0.1 STACK ;
  SAMENET M5  M5    0.1 STACK ;
  SAMENET M6  M6    0.1 STACK ;
  SAMENET V1  V1    0.1 ;
  SAMENET V2  V2    0.1 ;
  SAMENET V3  V3    0.1 ;
  SAMENET V4  V4    0.1 ;
  SAMENET V5  V5    0.1 ;
  SAMENET V1  V2    0.00 STACK ;
  SAMENET V2  V3    0.00 STACK ;
  SAMENET V3  V4    0.00 STACK ;
  SAMENET V4  V5    0.00 STACK ;
  SAMENET V1  V3    0.00 STACK ;
  SAMENET V2  V4    0.00 STACK ;
  SAMENET V3  V5    0.00 STACK ;
  SAMENET V1  V4    0.00 STACK ;
  SAMENET V2  V5    0.00 STACK ;
  SAMENET V1  V5    0.00 STACK ;
END SPACING


VIA via5 DEFAULT
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5

VIA via4 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4

VIA via3 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3

VIA via2 DEFAULT
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2

VIA via1 DEFAULT
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1


VIARULE via1Array GENERATE
  LAYER M1 ;
  DIRECTION HORIZONTAL ;
  OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via1Array


VIARULE via2Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via2Array


VIARULE via3Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via5Array

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
  LAYER M5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
END TURNM6


SITE  CoreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 4.71 ;
END  CoreSite

SITE  TDCoverSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  TDCoverSite

SITE  SBlockSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  SBlockSite

SITE  PortCellSite
    CLASS       PAD ;
    SIZE        0.0500 BY 0.0500 ;
END  PortCellSite

SITE  Core
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 4.71 ;
END  Core




MACRO AOI21
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN AOI21 0 -2.033 ;
  SIZE 2.08 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 -0.179 1 0.121 ;
      LAYER M2 ;
        RECT 0.86 -0.24 1 0.14 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 -0.179 1.512 0.121 ;
      LAYER M2 ;
        RECT 1.372 -0.24 1.512 0.14 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.655 -0.179 1.795 0.121 ;
        RECT 1.68 -0.532 1.77 1.161 ;
        RECT 1.238 -0.532 1.77 -0.442 ;
        RECT 1.238 -1.142 1.328 -0.442 ;
      LAYER M2 ;
        RECT 1.655 -0.24 1.795 0.14 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.08 -1.898 ;
        RECT 1.683 -2.033 1.773 -0.622 ;
        RECT 0.361 -2.033 0.451 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.08 2.677 ;
        RECT 0.765 0.441 0.855 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.278 0.261 1.368 1.161 ;
      RECT 0.375 0.261 0.465 1.161 ;
      RECT 0.375 0.261 1.368 0.351 ;
  END
  
END AOI21

MACRO AOI22
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN AOI22 0 -2.033 ;
  SIZE 2.6 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 -0.179 1 0.121 ;
      LAYER M2 ;
        RECT 0.86 -0.24 1 0.14 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 -0.179 1.512 0.121 ;
      LAYER M2 ;
        RECT 1.372 -0.24 1.512 0.14 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.154 -0.179 2.294 0.121 ;
      LAYER M2 ;
        RECT 2.154 -0.24 2.294 0.14 ;
      LAYER V1 ;
        RECT 2.174 -0.05 2.274 0.05 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.643 -0.179 1.783 0.121 ;
        RECT 1.673 -0.532 1.763 1.161 ;
        RECT 1.265 -0.532 1.763 -0.442 ;
        RECT 1.265 -1.142 1.355 -0.442 ;
      LAYER M2 ;
        RECT 1.643 -0.24 1.783 0.14 ;
      LAYER V1 ;
        RECT 1.663 -0.05 1.763 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.6 -1.898 ;
        RECT 2.192 -2.033 2.282 -0.622 ;
        RECT 0.361 -2.033 0.451 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.6 2.677 ;
        RECT 0.854 0.441 0.944 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.292 1.993 2.307 2.083 ;
      RECT 2.217 0.441 2.307 2.083 ;
      RECT 1.292 0.258 1.382 2.083 ;
      RECT 0.369 0.258 0.459 1.161 ;
      RECT 0.369 0.258 1.382 0.348 ;
  END
  
END AOI22

MACRO DFF
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN DFF 0 -2.033 ;
  SIZE 5.46 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.355 -0.179 2.495 0.121 ;
      LAYER M2 ;
        RECT 2.355 -0.24 2.495 0.14 ;
      LAYER V1 ;
        RECT 2.375 -0.05 2.475 0.05 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.308 -0.179 0.448 0.121 ;
      LAYER M2 ;
        RECT 0.308 -0.24 0.448 0.14 ;
      LAYER V1 ;
        RECT 0.328 -0.05 0.428 0.05 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.224 -0.179 3.364 0.121 ;
        RECT 3.249 -1.142 3.339 1.13 ;
      LAYER M2 ;
        RECT 3.224 -0.24 3.364 0.14 ;
      LAYER V1 ;
        RECT 3.244 -0.05 3.344 0.05 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.314 -0.179 1.454 0.121 ;
      LAYER M2 ;
        RECT 1.314 -0.24 1.454 0.14 ;
      LAYER V1 ;
        RECT 1.334 -0.05 1.434 0.05 ;
    END
  END R
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 5.46 -1.898 ;
        RECT 5.225 -2.033 5.315 -0.622 ;
        RECT 4.639 -2.033 4.729 -0.622 ;
        RECT 3.671 -2.033 3.761 -0.622 ;
        RECT 2.62 -2.033 2.71 -0.622 ;
        RECT 1.869 -2.033 1.959 -0.622 ;
        RECT 1.344 -2.033 1.434 -0.622 ;
        RECT 0.338 -2.033 0.428 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 5.46 2.677 ;
        RECT 4.639 0.41 4.729 2.677 ;
        RECT 3.671 0.41 3.761 2.677 ;
        RECT 2.465 0.41 2.555 2.677 ;
        RECT 1.301 0.441 1.391 2.677 ;
        RECT 0.338 0.441 0.428 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 5.225 -0.532 5.315 1.13 ;
      RECT 4.524 0.177 5.315 0.317 ;
      RECT 4.963 -0.532 5.315 -0.442 ;
      RECT 4.963 -1.142 5.053 -0.442 ;
      RECT 4.125 -1.142 4.215 1.13 ;
      RECT 3.556 0.177 4.215 0.317 ;
      RECT 4.125 -0.141 5.108 -0.001 ;
      RECT 2.881 1.256 3.327 1.346 ;
      RECT 2.882 -1.791 2.972 1.346 ;
      RECT 2.882 -1.756 3.569 -1.666 ;
      RECT 2.12 0.23 2.21 2.26 ;
      RECT 1.485 2.135 2.37 2.225 ;
      RECT 2.12 0.23 2.765 0.32 ;
      RECT 2.625 -0.532 2.765 0.32 ;
      RECT 2.12 -0.532 2.765 -0.442 ;
      RECT 2.12 -1.142 2.21 -0.442 ;
      RECT 1.869 0.031 1.959 1.561 ;
      RECT 1.191 0.211 1.959 0.351 ;
      RECT 1.606 0.031 1.959 0.121 ;
      RECT 1.606 -1.142 1.696 0.121 ;
      RECT 0.792 -1.526 0.882 1.161 ;
      RECT 0.792 -1.526 1.254 -1.436 ;
      RECT 3.857 2.367 4.534 2.457 ;
      RECT 2.65 1.436 3.577 1.526 ;
      RECT 2.65 1.902 3.577 1.992 ;
      RECT 2.65 2.135 3.577 2.225 ;
      RECT 2.9 2.368 3.577 2.458 ;
      RECT 2.65 1.669 3.123 1.759 ;
      RECT 2.049 -1.756 2.53 -1.666 ;
      RECT 1.49 1.669 2.03 1.759 ;
      RECT 1.485 1.902 1.971 1.992 ;
      RECT 0.737 -1.756 1.254 -1.666 ;
  END
  
END DFF

MACRO INVERTER
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN INVERTER 0 -2.033 ;
  SIZE 1.04 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.621 -0.179 0.761 0.121 ;
        RECT 0.646 -1.142 0.736 1.161 ;
      LAYER M2 ;
        RECT 0.621 -0.24 0.761 0.14 ;
      LAYER V1 ;
        RECT 0.641 -0.05 0.741 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 1.04 -1.898 ;
        RECT 0.341 -2.033 0.431 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 1.04 2.677 ;
        RECT 0.341 0.441 0.431 2.677 ;
    END
  END VDD!
  
END INVERTER

MACRO MUX21
  CLASS CORE ;
  ORIGIN 0 1.823 ;
  FOREIGN MUX21 0 -1.823 ;
  SIZE 3.12 BY 4.5 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.133 -0.107 1.319 0.121 ;
      LAYER M2 ;
        RECT 1.133 -0.14 1.319 0.14 ;
      LAYER V1 ;
        RECT 1.15 -0.05 1.25 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.156 -0.107 2.342 0.121 ;
      LAYER M2 ;
        RECT 2.156 -0.14 2.342 0.14 ;
      LAYER V1 ;
        RECT 2.173 -0.05 2.273 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.696 -0.107 2.882 0.121 ;
        RECT 2.705 -0.931 2.795 1.161 ;
      LAYER M2 ;
        RECT 2.696 -0.14 2.882 0.14 ;
      LAYER V1 ;
        RECT 2.696 -0.05 2.796 0.05 ;
    END
  END OUT
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.621 -0.107 0.807 0.121 ;
      LAYER M2 ;
        RECT 0.621 -0.14 0.807 0.14 ;
      LAYER V1 ;
        RECT 0.638 -0.05 0.738 0.05 ;
    END
  END S
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -1.823 3.12 -1.688 ;
        RECT 2.282 -1.823 2.372 -0.411 ;
        RECT 0.754 -1.823 0.844 -0.411 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 3.12 2.677 ;
        RECT 2.276 0.441 2.366 2.677 ;
        RECT 0.856 0.441 0.946 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.698 -1.515 1.788 1.161 ;
      RECT 0.369 -1.433 0.459 2.062 ;
  END
  
END MUX21

MACRO NAND2
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN NAND2 0 -2.033 ;
  SIZE 1.56 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.799 -0.179 0.939 0.121 ;
      LAYER M2 ;
        RECT 0.799 -0.24 0.939 0.14 ;
      LAYER V1 ;
        RECT 0.819 -0.05 0.919 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.082 -0.179 1.222 0.121 ;
        RECT 1.103 -1.142 1.193 1.131 ;
        RECT 0.341 0.211 1.193 0.301 ;
        RECT 0.341 0.211 0.431 1.131 ;
      LAYER M2 ;
        RECT 1.082 -0.24 1.222 0.14 ;
      LAYER V1 ;
        RECT 1.102 -0.05 1.202 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 1.56 -1.898 ;
        RECT 0.341 -2.033 0.431 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 1.56 2.677 ;
        RECT 0.725 0.411 0.815 2.677 ;
    END
  END VDD!
  
END NAND2

MACRO NAND3
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN NAND3 0 -2.033 ;
  SIZE 2.08 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 -0.179 1.512 0.121 ;
      LAYER M2 ;
        RECT 1.372 -0.24 1.512 0.14 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 -0.179 1 0.121 ;
      LAYER M2 ;
        RECT 0.86 -0.24 1 0.14 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.655 -0.179 1.795 0.121 ;
        RECT 1.679 -1.142 1.769 1.161 ;
        RECT 0.85 0.211 1.769 0.301 ;
        RECT 0.85 0.211 0.94 1.161 ;
      LAYER M2 ;
        RECT 1.655 -0.24 1.795 0.14 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.08 -1.898 ;
        RECT 0.377 -2.033 0.467 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.08 2.677 ;
        RECT 1.239 0.441 1.329 2.677 ;
        RECT 0.369 0.441 0.459 2.677 ;
    END
  END VDD!
  
END NAND3

MACRO NAND4
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN NAND4 0 -2.033 ;
  SIZE 2.6 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.884 -0.179 2.024 0.121 ;
      LAYER M2 ;
        RECT 1.884 -0.24 2.024 0.14 ;
      LAYER V1 ;
        RECT 1.904 -0.05 2.004 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 -0.179 1.512 0.121 ;
      LAYER M2 ;
        RECT 1.372 -0.24 1.512 0.14 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 -0.179 1 0.121 ;
      LAYER M2 ;
        RECT 0.86 -0.24 1 0.14 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.167 -0.179 2.307 0.121 ;
        RECT 0.854 0.211 2.282 0.301 ;
        RECT 2.192 -1.142 2.282 0.301 ;
        RECT 1.747 0.211 1.837 1.161 ;
        RECT 0.854 0.211 0.944 1.161 ;
      LAYER M2 ;
        RECT 2.167 -0.24 2.307 0.14 ;
      LAYER V1 ;
        RECT 2.187 -0.05 2.287 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.6 -1.898 ;
        RECT 0.377 -2.033 0.467 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.6 2.677 ;
        RECT 2.212 0.441 2.302 2.677 ;
        RECT 1.365 0.441 1.455 2.677 ;
        RECT 0.369 0.441 0.459 2.677 ;
    END
  END VDD!
  
END NAND4

MACRO NOR2
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN NOR2 0 -2.033 ;
  SIZE 1.56 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.799 -0.179 0.939 0.121 ;
      LAYER M2 ;
        RECT 0.799 -0.24 0.939 0.14 ;
      LAYER V1 ;
        RECT 0.819 -0.05 0.919 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.084 -0.179 1.224 0.121 ;
        RECT 1.102 -1.142 1.192 1.161 ;
        RECT 0.341 -0.532 1.192 -0.442 ;
        RECT 0.341 -1.142 0.431 -0.442 ;
      LAYER M2 ;
        RECT 1.084 -0.24 1.224 0.14 ;
      LAYER V1 ;
        RECT 1.102 -0.05 1.202 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 1.56 -1.898 ;
        RECT 0.726 -2.033 0.816 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 1.56 2.677 ;
        RECT 0.341 0.441 0.431 2.677 ;
    END
  END VDD!
  
END NOR2

MACRO NOR3
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN NOR3 0 -2.033 ;
  SIZE 2.08 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 -0.179 1 0.121 ;
      LAYER M2 ;
        RECT 0.86 -0.24 1 0.14 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 -0.179 1.512 0.121 ;
      LAYER M2 ;
        RECT 1.372 -0.24 1.512 0.14 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.655 -0.179 1.795 0.121 ;
        RECT 1.68 -1.142 1.77 1.161 ;
        RECT 0.856 -0.532 1.77 -0.442 ;
        RECT 0.856 -1.139 0.946 -0.442 ;
      LAYER M2 ;
        RECT 1.655 -0.24 1.795 0.14 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.08 -1.898 ;
        RECT 1.24 -2.033 1.33 -0.622 ;
        RECT 0.377 -2.033 0.467 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.08 2.677 ;
        RECT 0.369 0.441 0.459 2.677 ;
    END
  END VDD!
  
END NOR3

MACRO OAI21
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN OAI21 0 -2.033 ;
  SIZE 2.08 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 -0.179 1 0.121 ;
      LAYER M2 ;
        RECT 0.86 -0.24 1 0.14 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 -0.179 1.512 0.121 ;
      LAYER M2 ;
        RECT 1.372 -0.24 1.512 0.14 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.655 -0.107 1.795 0.121 ;
        RECT 1.269 0.211 1.77 0.301 ;
        RECT 1.68 -1.142 1.77 0.301 ;
        RECT 1.269 0.211 1.359 1.161 ;
      LAYER M2 ;
        RECT 1.655 -0.24 1.795 0.14 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.08 -1.898 ;
        RECT 0.854 -2.033 0.944 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.08 2.677 ;
        RECT 1.701 0.441 1.791 2.677 ;
        RECT 0.369 0.441 0.459 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 0.377 -0.532 1.329 -0.442 ;
      RECT 1.239 -1.142 1.329 -0.442 ;
      RECT 0.377 -1.142 0.467 -0.442 ;
  END
  
END OAI21

MACRO OAI22
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN OAI22 0 -2.033 ;
  SIZE 2.6 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.154 -0.179 2.294 0.121 ;
      LAYER M2 ;
        RECT 2.154 -0.24 2.294 0.14 ;
      LAYER V1 ;
        RECT 2.174 -0.05 2.274 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 -0.179 1.512 0.121 ;
      LAYER M2 ;
        RECT 1.372 -0.24 1.512 0.14 ;
      LAYER V1 ;
        RECT 1.392 -0.05 1.492 0.05 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 -0.179 1 0.121 ;
      LAYER M2 ;
        RECT 0.86 -0.24 1 0.14 ;
      LAYER V1 ;
        RECT 0.88 -0.05 0.98 0.05 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.657 -0.179 1.797 0.121 ;
        RECT 1.289 0.211 1.773 0.301 ;
        RECT 1.683 -1.142 1.773 0.301 ;
        RECT 1.289 0.211 1.379 1.161 ;
      LAYER M2 ;
        RECT 1.657 -0.24 1.797 0.14 ;
      LAYER V1 ;
        RECT 1.677 -0.05 1.777 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.6 -1.898 ;
        RECT 0.765 -2.033 0.855 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.6 2.677 ;
        RECT 2.218 0.441 2.308 2.677 ;
        RECT 0.369 0.441 0.459 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 0.377 -0.532 1.363 -0.442 ;
      RECT 1.273 -1.447 1.363 -0.442 ;
      RECT 0.377 -1.142 0.467 -0.442 ;
      RECT 2.191 -1.447 2.281 -0.622 ;
      RECT 1.273 -1.447 2.281 -1.357 ;
  END
  
END OAI22

MACRO TRI_INV
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN TRI_INV 0 -2.033 ;
  SIZE 2.34 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.618 -0.179 0.758 0.121 ;
      LAYER M2 ;
        RECT 0.618 -0.24 0.758 0.14 ;
      LAYER V1 ;
        RECT 0.638 -0.05 0.738 0.05 ;
    END
  END EN
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.13 -0.179 1.27 0.121 ;
      LAYER M2 ;
        RECT 1.13 -0.24 1.27 0.14 ;
      LAYER V1 ;
        RECT 1.15 -0.05 1.25 0.05 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.655 -0.179 1.795 0.121 ;
        RECT 1.68 -1.142 1.77 1.161 ;
      LAYER M2 ;
        RECT 1.655 -0.24 1.795 0.14 ;
      LAYER V1 ;
        RECT 1.675 -0.05 1.775 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 2.34 -1.898 ;
        RECT 0.751 -2.033 0.841 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 2.34 2.677 ;
        RECT 0.857 0.441 0.947 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.239 1.251 2.122 1.341 ;
      RECT 2.032 -1.637 2.122 1.341 ;
      RECT 1.239 0.441 1.329 1.341 ;
      RECT 1.241 -1.637 1.331 -0.622 ;
      RECT 1.241 -1.637 2.122 -1.547 ;
      RECT 0.275 -1.142 0.365 2.032 ;
  END
  
END TRI_INV

MACRO XOR2
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN XOR2 0 -2.033 ;
  SIZE 3.12 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.799 -0.179 0.939 0.121 ;
      LAYER M2 ;
        RECT 0.799 -0.24 0.939 0.14 ;
      LAYER V1 ;
        RECT 0.819 -0.05 0.919 0.05 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 -0.179 0.488 0.121 ;
      LAYER M2 ;
        RECT 0.348 -0.24 0.488 0.14 ;
      LAYER V1 ;
        RECT 0.368 -0.05 0.468 0.05 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.165 -0.179 2.305 0.121 ;
        RECT 2.188 -0.532 2.278 1.161 ;
        RECT 1.769 -0.532 2.278 -0.442 ;
        RECT 1.769 -1.142 1.859 -0.442 ;
      LAYER M2 ;
        RECT 2.165 -0.24 2.305 0.14 ;
      LAYER V1 ;
        RECT 2.185 -0.05 2.285 0.05 ;
    END
  END OUT
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -2.033 3.12 -1.898 ;
        RECT 2.683 -2.033 2.773 -0.622 ;
        RECT 1.369 -2.033 1.459 -0.622 ;
        RECT 0.341 -2.033 0.431 -0.622 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 2.549 3.12 2.677 ;
        RECT 1.248 0.441 1.338 2.677 ;
    END
  END VDD!
  OBS
    LAYER M1 ;
      RECT 1.762 1.251 2.785 1.341 ;
      RECT 2.695 0.441 2.785 1.341 ;
      RECT 1.762 0.441 1.852 1.341 ;
      RECT 0.341 0.211 0.431 1.161 ;
      RECT 0.341 0.211 1.455 0.301 ;
      RECT 1.365 -0.532 1.455 0.301 ;
      RECT 0.727 -0.532 1.455 -0.442 ;
      RECT 0.727 -1.142 0.817 -0.442 ;
  END
  
END XOR2

MACRO filler
  CLASS CORE ;
  ORIGIN 0 2.033 ;
  FOREIGN filler 0 -2.033 ;
  SIZE 0.26 BY 4.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN GND!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.076 -2.033 0.325 -1.898 ;
    END
  END GND!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.076 2.549 0.325 2.677 ;
    END
  END VDD!
  
END filler

END LIBRARY
