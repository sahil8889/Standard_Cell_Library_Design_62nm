// Created by ihdl
module matrix_vector_mult (
	clk, 
	rst_n, 
	matrix00, 
	matrix01, 
	matrix02, 
	matrix10, 
	matrix11, 
	matrix12, 
	matrix20, 
	matrix21, 
	matrix22, 
	vector_0, 
	vector_1, 
	vector_2, 
	result_0, 
	result_1, 
	result_2);
   input clk;
   input rst_n;
   input [7:0] matrix00;
   input [7:0] matrix01;
   input [7:0] matrix02;
   input [7:0] matrix10;
   input [7:0] matrix11;
   input [7:0] matrix12;
   input [7:0] matrix20;
   input [7:0] matrix21;
   input [7:0] matrix22;
   input [7:0] vector_0;
   input [7:0] vector_1;
   input [7:0] vector_2;
   output [15:0] result_0;
   output [15:0] result_1;
   output [15:0] result_2;

   // Internal wires
   wire N0;
   wire N1;
   wire N3;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N49;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N67;
   wire N68;
   wire N69;
   wire N70;
   wire N71;
   wire N72;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N129;
   wire N131;
   wire N132;
   wire N133;
   wire N134;
   wire N135;
   wire N136;
   wire N137;
   wire N138;
   wire N139;
   wire N140;
   wire N141;
   wire N142;
   wire N143;
   wire N144;
   wire N145;
   wire N146;
   wire N147;
   wire N148;
   wire N149;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N209;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire n1;
   wire \mult_21_3/FS_1/C[1][2][0] ;
   wire \mult_21_3/FS_1/C[1][2][1] ;
   wire \mult_21_3/FS_1/C[1][2][2] ;
   wire \mult_21_3/FS_1/C[1][2][3] ;
   wire \mult_21_3/FS_1/C[1][3][0] ;
   wire \mult_21_3/FS_1/C[1][3][1] ;
   wire \mult_21_3/FS_1/P[0][0][1] ;
   wire \mult_21_3/FS_1/P[0][0][2] ;
   wire \mult_21_3/FS_1/P[0][0][3] ;
   wire \mult_21_3/FS_1/P[0][1][1] ;
   wire \mult_21_3/FS_1/P[0][1][2] ;
   wire \mult_21_3/FS_1/P[0][1][3] ;
   wire \mult_21_3/FS_1/P[0][2][1] ;
   wire \mult_21_3/FS_1/P[0][2][2] ;
   wire \mult_21_3/FS_1/P[0][2][3] ;
   wire \mult_21_3/FS_1/P[0][3][1] ;
   wire \mult_21_3/FS_1/TEMP_P[0][0][0] ;
   wire \mult_21_3/FS_1/TEMP_P[0][1][0] ;
   wire \mult_21_3/FS_1/TEMP_P[0][2][0] ;
   wire \mult_21_3/FS_1/TEMP_P[0][2][1] ;
   wire \mult_21_3/FS_1/TEMP_P[0][2][2] ;
   wire \mult_21_3/FS_1/TEMP_P[0][3][0] ;
   wire \mult_21_3/FS_1/G[1][0][1] ;
   wire \mult_21_3/FS_1/G[1][0][2] ;
   wire \mult_21_3/FS_1/TEMP_G[0][2][1] ;
   wire \mult_21_3/FS_1/TEMP_G[0][2][2] ;
   wire \mult_21_3/FS_1/G_n_int[0][1][3] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][0] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][1] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][2] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][3] ;
   wire \mult_21_3/FS_1/G_n_int[0][3][0] ;
   wire \mult_21_3/FS_1/PG_int[0][2][0] ;
   wire \mult_21_3/FS_1/PG_int[0][2][1] ;
   wire \mult_21_3/FS_1/PG_int[0][2][2] ;
   wire \mult_21_3/FS_1/PG_int[0][2][3] ;
   wire \mult_21_3/FS_1/PG_int[0][3][0] ;
   wire \mult_21_3/FS_1/PG_int[0][3][1] ;
   wire \mult_21_3/A2[7] ;
   wire \mult_21_3/A2[8] ;
   wire \mult_21_3/A2[9] ;
   wire \mult_21_3/A2[10] ;
   wire \mult_21_3/A2[11] ;
   wire \mult_21_3/A2[12] ;
   wire \mult_21_3/A2[13] ;
   wire \mult_21_3/A1[0] ;
   wire \mult_21_3/A1[1] ;
   wire \mult_21_3/A1[2] ;
   wire \mult_21_3/A1[3] ;
   wire \mult_21_3/A1[4] ;
   wire \mult_21_3/A1[5] ;
   wire \mult_21_3/A1[6] ;
   wire \mult_21_3/A1[7] ;
   wire \mult_21_3/A1[8] ;
   wire \mult_21_3/A1[9] ;
   wire \mult_21_3/A1[10] ;
   wire \mult_21_3/A1[11] ;
   wire \mult_21_3/A1[12] ;
   wire \mult_21_3/ab[0][1] ;
   wire \mult_21_3/ab[0][2] ;
   wire \mult_21_3/ab[0][3] ;
   wire \mult_21_3/ab[0][4] ;
   wire \mult_21_3/ab[0][5] ;
   wire \mult_21_3/ab[0][6] ;
   wire \mult_21_3/ab[0][7] ;
   wire \mult_21_3/ab[1][0] ;
   wire \mult_21_3/ab[1][1] ;
   wire \mult_21_3/ab[1][2] ;
   wire \mult_21_3/ab[1][3] ;
   wire \mult_21_3/ab[1][4] ;
   wire \mult_21_3/ab[1][5] ;
   wire \mult_21_3/ab[1][6] ;
   wire \mult_21_3/ab[1][7] ;
   wire \mult_21_3/ab[2][0] ;
   wire \mult_21_3/ab[2][1] ;
   wire \mult_21_3/ab[2][2] ;
   wire \mult_21_3/ab[2][3] ;
   wire \mult_21_3/ab[2][4] ;
   wire \mult_21_3/ab[2][5] ;
   wire \mult_21_3/ab[2][6] ;
   wire \mult_21_3/ab[2][7] ;
   wire \mult_21_3/ab[3][0] ;
   wire \mult_21_3/ab[3][1] ;
   wire \mult_21_3/ab[3][2] ;
   wire \mult_21_3/ab[3][3] ;
   wire \mult_21_3/ab[3][4] ;
   wire \mult_21_3/ab[3][5] ;
   wire \mult_21_3/ab[3][6] ;
   wire \mult_21_3/ab[3][7] ;
   wire \mult_21_3/ab[4][0] ;
   wire \mult_21_3/ab[4][1] ;
   wire \mult_21_3/ab[4][2] ;
   wire \mult_21_3/ab[4][3] ;
   wire \mult_21_3/ab[4][4] ;
   wire \mult_21_3/ab[4][5] ;
   wire \mult_21_3/ab[4][6] ;
   wire \mult_21_3/ab[4][7] ;
   wire \mult_21_3/ab[5][0] ;
   wire \mult_21_3/ab[5][1] ;
   wire \mult_21_3/ab[5][2] ;
   wire \mult_21_3/ab[5][3] ;
   wire \mult_21_3/ab[5][4] ;
   wire \mult_21_3/ab[5][5] ;
   wire \mult_21_3/ab[5][6] ;
   wire \mult_21_3/ab[5][7] ;
   wire \mult_21_3/ab[6][0] ;
   wire \mult_21_3/ab[6][1] ;
   wire \mult_21_3/ab[6][2] ;
   wire \mult_21_3/ab[6][3] ;
   wire \mult_21_3/ab[6][4] ;
   wire \mult_21_3/ab[6][5] ;
   wire \mult_21_3/ab[6][6] ;
   wire \mult_21_3/ab[6][7] ;
   wire \mult_21_3/ab[7][0] ;
   wire \mult_21_3/ab[7][1] ;
   wire \mult_21_3/ab[7][2] ;
   wire \mult_21_3/ab[7][3] ;
   wire \mult_21_3/ab[7][4] ;
   wire \mult_21_3/ab[7][5] ;
   wire \mult_21_3/ab[7][6] ;
   wire \mult_21_3/ab[7][7] ;
   wire \mult_21_3/B_not[7] ;
   wire \mult_21_3/A_not[7] ;
   wire \mult_21_2/FS_1/C[1][2][0] ;
   wire \mult_21_2/FS_1/C[1][2][1] ;
   wire \mult_21_2/FS_1/C[1][2][2] ;
   wire \mult_21_2/FS_1/C[1][2][3] ;
   wire \mult_21_2/FS_1/C[1][3][0] ;
   wire \mult_21_2/FS_1/C[1][3][1] ;
   wire \mult_21_2/FS_1/P[0][0][1] ;
   wire \mult_21_2/FS_1/P[0][0][2] ;
   wire \mult_21_2/FS_1/P[0][0][3] ;
   wire \mult_21_2/FS_1/P[0][1][1] ;
   wire \mult_21_2/FS_1/P[0][1][2] ;
   wire \mult_21_2/FS_1/P[0][1][3] ;
   wire \mult_21_2/FS_1/P[0][2][1] ;
   wire \mult_21_2/FS_1/P[0][2][2] ;
   wire \mult_21_2/FS_1/P[0][2][3] ;
   wire \mult_21_2/FS_1/P[0][3][1] ;
   wire \mult_21_2/FS_1/TEMP_P[0][0][0] ;
   wire \mult_21_2/FS_1/TEMP_P[0][1][0] ;
   wire \mult_21_2/FS_1/TEMP_P[0][2][0] ;
   wire \mult_21_2/FS_1/TEMP_P[0][2][1] ;
   wire \mult_21_2/FS_1/TEMP_P[0][2][2] ;
   wire \mult_21_2/FS_1/TEMP_P[0][3][0] ;
   wire \mult_21_2/FS_1/G[1][0][1] ;
   wire \mult_21_2/FS_1/G[1][0][2] ;
   wire \mult_21_2/FS_1/TEMP_G[0][2][1] ;
   wire \mult_21_2/FS_1/TEMP_G[0][2][2] ;
   wire \mult_21_2/FS_1/G_n_int[0][1][3] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][0] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][1] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][2] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][3] ;
   wire \mult_21_2/FS_1/G_n_int[0][3][0] ;
   wire \mult_21_2/FS_1/PG_int[0][2][0] ;
   wire \mult_21_2/FS_1/PG_int[0][2][1] ;
   wire \mult_21_2/FS_1/PG_int[0][2][2] ;
   wire \mult_21_2/FS_1/PG_int[0][2][3] ;
   wire \mult_21_2/FS_1/PG_int[0][3][0] ;
   wire \mult_21_2/FS_1/PG_int[0][3][1] ;
   wire \mult_21_2/A2[7] ;
   wire \mult_21_2/A2[8] ;
   wire \mult_21_2/A2[9] ;
   wire \mult_21_2/A2[10] ;
   wire \mult_21_2/A2[11] ;
   wire \mult_21_2/A2[12] ;
   wire \mult_21_2/A2[13] ;
   wire \mult_21_2/A1[0] ;
   wire \mult_21_2/A1[1] ;
   wire \mult_21_2/A1[2] ;
   wire \mult_21_2/A1[3] ;
   wire \mult_21_2/A1[4] ;
   wire \mult_21_2/A1[5] ;
   wire \mult_21_2/A1[6] ;
   wire \mult_21_2/A1[7] ;
   wire \mult_21_2/A1[8] ;
   wire \mult_21_2/A1[9] ;
   wire \mult_21_2/A1[10] ;
   wire \mult_21_2/A1[11] ;
   wire \mult_21_2/A1[12] ;
   wire \mult_21_2/ab[0][1] ;
   wire \mult_21_2/ab[0][2] ;
   wire \mult_21_2/ab[0][3] ;
   wire \mult_21_2/ab[0][4] ;
   wire \mult_21_2/ab[0][5] ;
   wire \mult_21_2/ab[0][6] ;
   wire \mult_21_2/ab[0][7] ;
   wire \mult_21_2/ab[1][0] ;
   wire \mult_21_2/ab[1][1] ;
   wire \mult_21_2/ab[1][2] ;
   wire \mult_21_2/ab[1][3] ;
   wire \mult_21_2/ab[1][4] ;
   wire \mult_21_2/ab[1][5] ;
   wire \mult_21_2/ab[1][6] ;
   wire \mult_21_2/ab[1][7] ;
   wire \mult_21_2/ab[2][0] ;
   wire \mult_21_2/ab[2][1] ;
   wire \mult_21_2/ab[2][2] ;
   wire \mult_21_2/ab[2][3] ;
   wire \mult_21_2/ab[2][4] ;
   wire \mult_21_2/ab[2][5] ;
   wire \mult_21_2/ab[2][6] ;
   wire \mult_21_2/ab[2][7] ;
   wire \mult_21_2/ab[3][0] ;
   wire \mult_21_2/ab[3][1] ;
   wire \mult_21_2/ab[3][2] ;
   wire \mult_21_2/ab[3][3] ;
   wire \mult_21_2/ab[3][4] ;
   wire \mult_21_2/ab[3][5] ;
   wire \mult_21_2/ab[3][6] ;
   wire \mult_21_2/ab[3][7] ;
   wire \mult_21_2/ab[4][0] ;
   wire \mult_21_2/ab[4][1] ;
   wire \mult_21_2/ab[4][2] ;
   wire \mult_21_2/ab[4][3] ;
   wire \mult_21_2/ab[4][4] ;
   wire \mult_21_2/ab[4][5] ;
   wire \mult_21_2/ab[4][6] ;
   wire \mult_21_2/ab[4][7] ;
   wire \mult_21_2/ab[5][0] ;
   wire \mult_21_2/ab[5][1] ;
   wire \mult_21_2/ab[5][2] ;
   wire \mult_21_2/ab[5][3] ;
   wire \mult_21_2/ab[5][4] ;
   wire \mult_21_2/ab[5][5] ;
   wire \mult_21_2/ab[5][6] ;
   wire \mult_21_2/ab[5][7] ;
   wire \mult_21_2/ab[6][0] ;
   wire \mult_21_2/ab[6][1] ;
   wire \mult_21_2/ab[6][2] ;
   wire \mult_21_2/ab[6][3] ;
   wire \mult_21_2/ab[6][4] ;
   wire \mult_21_2/ab[6][5] ;
   wire \mult_21_2/ab[6][6] ;
   wire \mult_21_2/ab[6][7] ;
   wire \mult_21_2/ab[7][0] ;
   wire \mult_21_2/ab[7][1] ;
   wire \mult_21_2/ab[7][2] ;
   wire \mult_21_2/ab[7][3] ;
   wire \mult_21_2/ab[7][4] ;
   wire \mult_21_2/ab[7][5] ;
   wire \mult_21_2/ab[7][6] ;
   wire \mult_21_2/ab[7][7] ;
   wire \mult_21_2/B_not[7] ;
   wire \mult_21_2/A_not[7] ;
   wire \mult_21/FS_1/C[1][2][0] ;
   wire \mult_21/FS_1/C[1][2][1] ;
   wire \mult_21/FS_1/C[1][2][2] ;
   wire \mult_21/FS_1/C[1][2][3] ;
   wire \mult_21/FS_1/C[1][3][0] ;
   wire \mult_21/FS_1/C[1][3][1] ;
   wire \mult_21/FS_1/P[0][0][1] ;
   wire \mult_21/FS_1/P[0][0][2] ;
   wire \mult_21/FS_1/P[0][0][3] ;
   wire \mult_21/FS_1/P[0][1][1] ;
   wire \mult_21/FS_1/P[0][1][2] ;
   wire \mult_21/FS_1/P[0][1][3] ;
   wire \mult_21/FS_1/P[0][2][1] ;
   wire \mult_21/FS_1/P[0][2][2] ;
   wire \mult_21/FS_1/P[0][2][3] ;
   wire \mult_21/FS_1/P[0][3][1] ;
   wire \mult_21/FS_1/TEMP_P[0][0][0] ;
   wire \mult_21/FS_1/TEMP_P[0][1][0] ;
   wire \mult_21/FS_1/TEMP_P[0][2][0] ;
   wire \mult_21/FS_1/TEMP_P[0][2][1] ;
   wire \mult_21/FS_1/TEMP_P[0][2][2] ;
   wire \mult_21/FS_1/TEMP_P[0][3][0] ;
   wire \mult_21/FS_1/G[1][0][1] ;
   wire \mult_21/FS_1/G[1][0][2] ;
   wire \mult_21/FS_1/TEMP_G[0][2][1] ;
   wire \mult_21/FS_1/TEMP_G[0][2][2] ;
   wire \mult_21/FS_1/G_n_int[0][1][3] ;
   wire \mult_21/FS_1/G_n_int[0][2][0] ;
   wire \mult_21/FS_1/G_n_int[0][2][1] ;
   wire \mult_21/FS_1/G_n_int[0][2][2] ;
   wire \mult_21/FS_1/G_n_int[0][2][3] ;
   wire \mult_21/FS_1/G_n_int[0][3][0] ;
   wire \mult_21/FS_1/PG_int[0][2][0] ;
   wire \mult_21/FS_1/PG_int[0][2][1] ;
   wire \mult_21/FS_1/PG_int[0][2][2] ;
   wire \mult_21/FS_1/PG_int[0][2][3] ;
   wire \mult_21/FS_1/PG_int[0][3][0] ;
   wire \mult_21/FS_1/PG_int[0][3][1] ;
   wire \mult_21/A2[7] ;
   wire \mult_21/A2[8] ;
   wire \mult_21/A2[9] ;
   wire \mult_21/A2[10] ;
   wire \mult_21/A2[11] ;
   wire \mult_21/A2[12] ;
   wire \mult_21/A2[13] ;
   wire \mult_21/A1[0] ;
   wire \mult_21/A1[1] ;
   wire \mult_21/A1[2] ;
   wire \mult_21/A1[3] ;
   wire \mult_21/A1[4] ;
   wire \mult_21/A1[5] ;
   wire \mult_21/A1[6] ;
   wire \mult_21/A1[7] ;
   wire \mult_21/A1[8] ;
   wire \mult_21/A1[9] ;
   wire \mult_21/A1[10] ;
   wire \mult_21/A1[11] ;
   wire \mult_21/A1[12] ;
   wire \mult_21/ab[0][1] ;
   wire \mult_21/ab[0][2] ;
   wire \mult_21/ab[0][3] ;
   wire \mult_21/ab[0][4] ;
   wire \mult_21/ab[0][5] ;
   wire \mult_21/ab[0][6] ;
   wire \mult_21/ab[0][7] ;
   wire \mult_21/ab[1][0] ;
   wire \mult_21/ab[1][1] ;
   wire \mult_21/ab[1][2] ;
   wire \mult_21/ab[1][3] ;
   wire \mult_21/ab[1][4] ;
   wire \mult_21/ab[1][5] ;
   wire \mult_21/ab[1][6] ;
   wire \mult_21/ab[1][7] ;
   wire \mult_21/ab[2][0] ;
   wire \mult_21/ab[2][1] ;
   wire \mult_21/ab[2][2] ;
   wire \mult_21/ab[2][3] ;
   wire \mult_21/ab[2][4] ;
   wire \mult_21/ab[2][5] ;
   wire \mult_21/ab[2][6] ;
   wire \mult_21/ab[2][7] ;
   wire \mult_21/ab[3][0] ;
   wire \mult_21/ab[3][1] ;
   wire \mult_21/ab[3][2] ;
   wire \mult_21/ab[3][3] ;
   wire \mult_21/ab[3][4] ;
   wire \mult_21/ab[3][5] ;
   wire \mult_21/ab[3][6] ;
   wire \mult_21/ab[3][7] ;
   wire \mult_21/ab[4][0] ;
   wire \mult_21/ab[4][1] ;
   wire \mult_21/ab[4][2] ;
   wire \mult_21/ab[4][3] ;
   wire \mult_21/ab[4][4] ;
   wire \mult_21/ab[4][5] ;
   wire \mult_21/ab[4][6] ;
   wire \mult_21/ab[4][7] ;
   wire \mult_21/ab[5][0] ;
   wire \mult_21/ab[5][1] ;
   wire \mult_21/ab[5][2] ;
   wire \mult_21/ab[5][3] ;
   wire \mult_21/ab[5][4] ;
   wire \mult_21/ab[5][5] ;
   wire \mult_21/ab[5][6] ;
   wire \mult_21/ab[5][7] ;
   wire \mult_21/ab[6][0] ;
   wire \mult_21/ab[6][1] ;
   wire \mult_21/ab[6][2] ;
   wire \mult_21/ab[6][3] ;
   wire \mult_21/ab[6][4] ;
   wire \mult_21/ab[6][5] ;
   wire \mult_21/ab[6][6] ;
   wire \mult_21/ab[6][7] ;
   wire \mult_21/ab[7][0] ;
   wire \mult_21/ab[7][1] ;
   wire \mult_21/ab[7][2] ;
   wire \mult_21/ab[7][3] ;
   wire \mult_21/ab[7][4] ;
   wire \mult_21/ab[7][5] ;
   wire \mult_21/ab[7][6] ;
   wire \mult_21/ab[7][7] ;
   wire \mult_21/B_not[7] ;
   wire \mult_21/A_not[7] ;
   wire \mult_20_3/FS_1/C[1][2][0] ;
   wire \mult_20_3/FS_1/C[1][2][1] ;
   wire \mult_20_3/FS_1/C[1][2][2] ;
   wire \mult_20_3/FS_1/C[1][2][3] ;
   wire \mult_20_3/FS_1/C[1][3][0] ;
   wire \mult_20_3/FS_1/C[1][3][1] ;
   wire \mult_20_3/FS_1/P[0][0][1] ;
   wire \mult_20_3/FS_1/P[0][0][2] ;
   wire \mult_20_3/FS_1/P[0][0][3] ;
   wire \mult_20_3/FS_1/P[0][1][1] ;
   wire \mult_20_3/FS_1/P[0][1][2] ;
   wire \mult_20_3/FS_1/P[0][1][3] ;
   wire \mult_20_3/FS_1/P[0][2][1] ;
   wire \mult_20_3/FS_1/P[0][2][2] ;
   wire \mult_20_3/FS_1/P[0][2][3] ;
   wire \mult_20_3/FS_1/P[0][3][1] ;
   wire \mult_20_3/FS_1/TEMP_P[0][0][0] ;
   wire \mult_20_3/FS_1/TEMP_P[0][1][0] ;
   wire \mult_20_3/FS_1/TEMP_P[0][2][0] ;
   wire \mult_20_3/FS_1/TEMP_P[0][2][1] ;
   wire \mult_20_3/FS_1/TEMP_P[0][2][2] ;
   wire \mult_20_3/FS_1/TEMP_P[0][3][0] ;
   wire \mult_20_3/FS_1/G[1][0][1] ;
   wire \mult_20_3/FS_1/G[1][0][2] ;
   wire \mult_20_3/FS_1/TEMP_G[0][2][1] ;
   wire \mult_20_3/FS_1/TEMP_G[0][2][2] ;
   wire \mult_20_3/FS_1/G_n_int[0][1][3] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][0] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][1] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][2] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][3] ;
   wire \mult_20_3/FS_1/G_n_int[0][3][0] ;
   wire \mult_20_3/FS_1/PG_int[0][2][0] ;
   wire \mult_20_3/FS_1/PG_int[0][2][1] ;
   wire \mult_20_3/FS_1/PG_int[0][2][2] ;
   wire \mult_20_3/FS_1/PG_int[0][2][3] ;
   wire \mult_20_3/FS_1/PG_int[0][3][0] ;
   wire \mult_20_3/FS_1/PG_int[0][3][1] ;
   wire \mult_20_3/A2[7] ;
   wire \mult_20_3/A2[8] ;
   wire \mult_20_3/A2[9] ;
   wire \mult_20_3/A2[10] ;
   wire \mult_20_3/A2[11] ;
   wire \mult_20_3/A2[12] ;
   wire \mult_20_3/A2[13] ;
   wire \mult_20_3/A1[0] ;
   wire \mult_20_3/A1[1] ;
   wire \mult_20_3/A1[2] ;
   wire \mult_20_3/A1[3] ;
   wire \mult_20_3/A1[4] ;
   wire \mult_20_3/A1[5] ;
   wire \mult_20_3/A1[6] ;
   wire \mult_20_3/A1[7] ;
   wire \mult_20_3/A1[8] ;
   wire \mult_20_3/A1[9] ;
   wire \mult_20_3/A1[10] ;
   wire \mult_20_3/A1[11] ;
   wire \mult_20_3/A1[12] ;
   wire \mult_20_3/ab[0][1] ;
   wire \mult_20_3/ab[0][2] ;
   wire \mult_20_3/ab[0][3] ;
   wire \mult_20_3/ab[0][4] ;
   wire \mult_20_3/ab[0][5] ;
   wire \mult_20_3/ab[0][6] ;
   wire \mult_20_3/ab[0][7] ;
   wire \mult_20_3/ab[1][0] ;
   wire \mult_20_3/ab[1][1] ;
   wire \mult_20_3/ab[1][2] ;
   wire \mult_20_3/ab[1][3] ;
   wire \mult_20_3/ab[1][4] ;
   wire \mult_20_3/ab[1][5] ;
   wire \mult_20_3/ab[1][6] ;
   wire \mult_20_3/ab[1][7] ;
   wire \mult_20_3/ab[2][0] ;
   wire \mult_20_3/ab[2][1] ;
   wire \mult_20_3/ab[2][2] ;
   wire \mult_20_3/ab[2][3] ;
   wire \mult_20_3/ab[2][4] ;
   wire \mult_20_3/ab[2][5] ;
   wire \mult_20_3/ab[2][6] ;
   wire \mult_20_3/ab[2][7] ;
   wire \mult_20_3/ab[3][0] ;
   wire \mult_20_3/ab[3][1] ;
   wire \mult_20_3/ab[3][2] ;
   wire \mult_20_3/ab[3][3] ;
   wire \mult_20_3/ab[3][4] ;
   wire \mult_20_3/ab[3][5] ;
   wire \mult_20_3/ab[3][6] ;
   wire \mult_20_3/ab[3][7] ;
   wire \mult_20_3/ab[4][0] ;
   wire \mult_20_3/ab[4][1] ;
   wire \mult_20_3/ab[4][2] ;
   wire \mult_20_3/ab[4][3] ;
   wire \mult_20_3/ab[4][4] ;
   wire \mult_20_3/ab[4][5] ;
   wire \mult_20_3/ab[4][6] ;
   wire \mult_20_3/ab[4][7] ;
   wire \mult_20_3/ab[5][0] ;
   wire \mult_20_3/ab[5][1] ;
   wire \mult_20_3/ab[5][2] ;
   wire \mult_20_3/ab[5][3] ;
   wire \mult_20_3/ab[5][4] ;
   wire \mult_20_3/ab[5][5] ;
   wire \mult_20_3/ab[5][6] ;
   wire \mult_20_3/ab[5][7] ;
   wire \mult_20_3/ab[6][0] ;
   wire \mult_20_3/ab[6][1] ;
   wire \mult_20_3/ab[6][2] ;
   wire \mult_20_3/ab[6][3] ;
   wire \mult_20_3/ab[6][4] ;
   wire \mult_20_3/ab[6][5] ;
   wire \mult_20_3/ab[6][6] ;
   wire \mult_20_3/ab[6][7] ;
   wire \mult_20_3/ab[7][0] ;
   wire \mult_20_3/ab[7][1] ;
   wire \mult_20_3/ab[7][2] ;
   wire \mult_20_3/ab[7][3] ;
   wire \mult_20_3/ab[7][4] ;
   wire \mult_20_3/ab[7][5] ;
   wire \mult_20_3/ab[7][6] ;
   wire \mult_20_3/ab[7][7] ;
   wire \mult_20_3/B_not[7] ;
   wire \mult_20_3/A_not[7] ;
   wire \mult_20_2/FS_1/C[1][2][0] ;
   wire \mult_20_2/FS_1/C[1][2][1] ;
   wire \mult_20_2/FS_1/C[1][2][2] ;
   wire \mult_20_2/FS_1/C[1][2][3] ;
   wire \mult_20_2/FS_1/C[1][3][0] ;
   wire \mult_20_2/FS_1/C[1][3][1] ;
   wire \mult_20_2/FS_1/P[0][0][1] ;
   wire \mult_20_2/FS_1/P[0][0][2] ;
   wire \mult_20_2/FS_1/P[0][0][3] ;
   wire \mult_20_2/FS_1/P[0][1][1] ;
   wire \mult_20_2/FS_1/P[0][1][2] ;
   wire \mult_20_2/FS_1/P[0][1][3] ;
   wire \mult_20_2/FS_1/P[0][2][1] ;
   wire \mult_20_2/FS_1/P[0][2][2] ;
   wire \mult_20_2/FS_1/P[0][2][3] ;
   wire \mult_20_2/FS_1/P[0][3][1] ;
   wire \mult_20_2/FS_1/TEMP_P[0][0][0] ;
   wire \mult_20_2/FS_1/TEMP_P[0][1][0] ;
   wire \mult_20_2/FS_1/TEMP_P[0][2][0] ;
   wire \mult_20_2/FS_1/TEMP_P[0][2][1] ;
   wire \mult_20_2/FS_1/TEMP_P[0][2][2] ;
   wire \mult_20_2/FS_1/TEMP_P[0][3][0] ;
   wire \mult_20_2/FS_1/G[1][0][1] ;
   wire \mult_20_2/FS_1/G[1][0][2] ;
   wire \mult_20_2/FS_1/TEMP_G[0][2][1] ;
   wire \mult_20_2/FS_1/TEMP_G[0][2][2] ;
   wire \mult_20_2/FS_1/G_n_int[0][1][3] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][0] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][1] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][2] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][3] ;
   wire \mult_20_2/FS_1/G_n_int[0][3][0] ;
   wire \mult_20_2/FS_1/PG_int[0][2][0] ;
   wire \mult_20_2/FS_1/PG_int[0][2][1] ;
   wire \mult_20_2/FS_1/PG_int[0][2][2] ;
   wire \mult_20_2/FS_1/PG_int[0][2][3] ;
   wire \mult_20_2/FS_1/PG_int[0][3][0] ;
   wire \mult_20_2/FS_1/PG_int[0][3][1] ;
   wire \mult_20_2/A2[7] ;
   wire \mult_20_2/A2[8] ;
   wire \mult_20_2/A2[9] ;
   wire \mult_20_2/A2[10] ;
   wire \mult_20_2/A2[11] ;
   wire \mult_20_2/A2[12] ;
   wire \mult_20_2/A2[13] ;
   wire \mult_20_2/A1[0] ;
   wire \mult_20_2/A1[1] ;
   wire \mult_20_2/A1[2] ;
   wire \mult_20_2/A1[3] ;
   wire \mult_20_2/A1[4] ;
   wire \mult_20_2/A1[5] ;
   wire \mult_20_2/A1[6] ;
   wire \mult_20_2/A1[7] ;
   wire \mult_20_2/A1[8] ;
   wire \mult_20_2/A1[9] ;
   wire \mult_20_2/A1[10] ;
   wire \mult_20_2/A1[11] ;
   wire \mult_20_2/A1[12] ;
   wire \mult_20_2/ab[0][1] ;
   wire \mult_20_2/ab[0][2] ;
   wire \mult_20_2/ab[0][3] ;
   wire \mult_20_2/ab[0][4] ;
   wire \mult_20_2/ab[0][5] ;
   wire \mult_20_2/ab[0][6] ;
   wire \mult_20_2/ab[0][7] ;
   wire \mult_20_2/ab[1][0] ;
   wire \mult_20_2/ab[1][1] ;
   wire \mult_20_2/ab[1][2] ;
   wire \mult_20_2/ab[1][3] ;
   wire \mult_20_2/ab[1][4] ;
   wire \mult_20_2/ab[1][5] ;
   wire \mult_20_2/ab[1][6] ;
   wire \mult_20_2/ab[1][7] ;
   wire \mult_20_2/ab[2][0] ;
   wire \mult_20_2/ab[2][1] ;
   wire \mult_20_2/ab[2][2] ;
   wire \mult_20_2/ab[2][3] ;
   wire \mult_20_2/ab[2][4] ;
   wire \mult_20_2/ab[2][5] ;
   wire \mult_20_2/ab[2][6] ;
   wire \mult_20_2/ab[2][7] ;
   wire \mult_20_2/ab[3][0] ;
   wire \mult_20_2/ab[3][1] ;
   wire \mult_20_2/ab[3][2] ;
   wire \mult_20_2/ab[3][3] ;
   wire \mult_20_2/ab[3][4] ;
   wire \mult_20_2/ab[3][5] ;
   wire \mult_20_2/ab[3][6] ;
   wire \mult_20_2/ab[3][7] ;
   wire \mult_20_2/ab[4][0] ;
   wire \mult_20_2/ab[4][1] ;
   wire \mult_20_2/ab[4][2] ;
   wire \mult_20_2/ab[4][3] ;
   wire \mult_20_2/ab[4][4] ;
   wire \mult_20_2/ab[4][5] ;
   wire \mult_20_2/ab[4][6] ;
   wire \mult_20_2/ab[4][7] ;
   wire \mult_20_2/ab[5][0] ;
   wire \mult_20_2/ab[5][1] ;
   wire \mult_20_2/ab[5][2] ;
   wire \mult_20_2/ab[5][3] ;
   wire \mult_20_2/ab[5][4] ;
   wire \mult_20_2/ab[5][5] ;
   wire \mult_20_2/ab[5][6] ;
   wire \mult_20_2/ab[5][7] ;
   wire \mult_20_2/ab[6][0] ;
   wire \mult_20_2/ab[6][1] ;
   wire \mult_20_2/ab[6][2] ;
   wire \mult_20_2/ab[6][3] ;
   wire \mult_20_2/ab[6][4] ;
   wire \mult_20_2/ab[6][5] ;
   wire \mult_20_2/ab[6][6] ;
   wire \mult_20_2/ab[6][7] ;
   wire \mult_20_2/ab[7][0] ;
   wire \mult_20_2/ab[7][1] ;
   wire \mult_20_2/ab[7][2] ;
   wire \mult_20_2/ab[7][3] ;
   wire \mult_20_2/ab[7][4] ;
   wire \mult_20_2/ab[7][5] ;
   wire \mult_20_2/ab[7][6] ;
   wire \mult_20_2/ab[7][7] ;
   wire \mult_20_2/B_not[7] ;
   wire \mult_20_2/A_not[7] ;
   wire \mult_20/FS_1/C[1][2][0] ;
   wire \mult_20/FS_1/C[1][2][1] ;
   wire \mult_20/FS_1/C[1][2][2] ;
   wire \mult_20/FS_1/C[1][2][3] ;
   wire \mult_20/FS_1/C[1][3][0] ;
   wire \mult_20/FS_1/C[1][3][1] ;
   wire \mult_20/FS_1/P[0][0][1] ;
   wire \mult_20/FS_1/P[0][0][2] ;
   wire \mult_20/FS_1/P[0][0][3] ;
   wire \mult_20/FS_1/P[0][1][1] ;
   wire \mult_20/FS_1/P[0][1][2] ;
   wire \mult_20/FS_1/P[0][1][3] ;
   wire \mult_20/FS_1/P[0][2][1] ;
   wire \mult_20/FS_1/P[0][2][2] ;
   wire \mult_20/FS_1/P[0][2][3] ;
   wire \mult_20/FS_1/P[0][3][1] ;
   wire \mult_20/FS_1/TEMP_P[0][0][0] ;
   wire \mult_20/FS_1/TEMP_P[0][1][0] ;
   wire \mult_20/FS_1/TEMP_P[0][2][0] ;
   wire \mult_20/FS_1/TEMP_P[0][2][1] ;
   wire \mult_20/FS_1/TEMP_P[0][2][2] ;
   wire \mult_20/FS_1/TEMP_P[0][3][0] ;
   wire \mult_20/FS_1/G[1][0][1] ;
   wire \mult_20/FS_1/G[1][0][2] ;
   wire \mult_20/FS_1/TEMP_G[0][2][1] ;
   wire \mult_20/FS_1/TEMP_G[0][2][2] ;
   wire \mult_20/FS_1/G_n_int[0][1][3] ;
   wire \mult_20/FS_1/G_n_int[0][2][0] ;
   wire \mult_20/FS_1/G_n_int[0][2][1] ;
   wire \mult_20/FS_1/G_n_int[0][2][2] ;
   wire \mult_20/FS_1/G_n_int[0][2][3] ;
   wire \mult_20/FS_1/G_n_int[0][3][0] ;
   wire \mult_20/FS_1/PG_int[0][2][0] ;
   wire \mult_20/FS_1/PG_int[0][2][1] ;
   wire \mult_20/FS_1/PG_int[0][2][2] ;
   wire \mult_20/FS_1/PG_int[0][2][3] ;
   wire \mult_20/FS_1/PG_int[0][3][0] ;
   wire \mult_20/FS_1/PG_int[0][3][1] ;
   wire \mult_20/A2[7] ;
   wire \mult_20/A2[8] ;
   wire \mult_20/A2[9] ;
   wire \mult_20/A2[10] ;
   wire \mult_20/A2[11] ;
   wire \mult_20/A2[12] ;
   wire \mult_20/A2[13] ;
   wire \mult_20/A1[0] ;
   wire \mult_20/A1[1] ;
   wire \mult_20/A1[2] ;
   wire \mult_20/A1[3] ;
   wire \mult_20/A1[4] ;
   wire \mult_20/A1[5] ;
   wire \mult_20/A1[6] ;
   wire \mult_20/A1[7] ;
   wire \mult_20/A1[8] ;
   wire \mult_20/A1[9] ;
   wire \mult_20/A1[10] ;
   wire \mult_20/A1[11] ;
   wire \mult_20/A1[12] ;
   wire \mult_20/ab[0][1] ;
   wire \mult_20/ab[0][2] ;
   wire \mult_20/ab[0][3] ;
   wire \mult_20/ab[0][4] ;
   wire \mult_20/ab[0][5] ;
   wire \mult_20/ab[0][6] ;
   wire \mult_20/ab[0][7] ;
   wire \mult_20/ab[1][0] ;
   wire \mult_20/ab[1][1] ;
   wire \mult_20/ab[1][2] ;
   wire \mult_20/ab[1][3] ;
   wire \mult_20/ab[1][4] ;
   wire \mult_20/ab[1][5] ;
   wire \mult_20/ab[1][6] ;
   wire \mult_20/ab[1][7] ;
   wire \mult_20/ab[2][0] ;
   wire \mult_20/ab[2][1] ;
   wire \mult_20/ab[2][2] ;
   wire \mult_20/ab[2][3] ;
   wire \mult_20/ab[2][4] ;
   wire \mult_20/ab[2][5] ;
   wire \mult_20/ab[2][6] ;
   wire \mult_20/ab[2][7] ;
   wire \mult_20/ab[3][0] ;
   wire \mult_20/ab[3][1] ;
   wire \mult_20/ab[3][2] ;
   wire \mult_20/ab[3][3] ;
   wire \mult_20/ab[3][4] ;
   wire \mult_20/ab[3][5] ;
   wire \mult_20/ab[3][6] ;
   wire \mult_20/ab[3][7] ;
   wire \mult_20/ab[4][0] ;
   wire \mult_20/ab[4][1] ;
   wire \mult_20/ab[4][2] ;
   wire \mult_20/ab[4][3] ;
   wire \mult_20/ab[4][4] ;
   wire \mult_20/ab[4][5] ;
   wire \mult_20/ab[4][6] ;
   wire \mult_20/ab[4][7] ;
   wire \mult_20/ab[5][0] ;
   wire \mult_20/ab[5][1] ;
   wire \mult_20/ab[5][2] ;
   wire \mult_20/ab[5][3] ;
   wire \mult_20/ab[5][4] ;
   wire \mult_20/ab[5][5] ;
   wire \mult_20/ab[5][6] ;
   wire \mult_20/ab[5][7] ;
   wire \mult_20/ab[6][0] ;
   wire \mult_20/ab[6][1] ;
   wire \mult_20/ab[6][2] ;
   wire \mult_20/ab[6][3] ;
   wire \mult_20/ab[6][4] ;
   wire \mult_20/ab[6][5] ;
   wire \mult_20/ab[6][6] ;
   wire \mult_20/ab[6][7] ;
   wire \mult_20/ab[7][0] ;
   wire \mult_20/ab[7][1] ;
   wire \mult_20/ab[7][2] ;
   wire \mult_20/ab[7][3] ;
   wire \mult_20/ab[7][4] ;
   wire \mult_20/ab[7][5] ;
   wire \mult_20/ab[7][6] ;
   wire \mult_20/ab[7][7] ;
   wire \mult_20/B_not[7] ;
   wire \mult_20/A_not[7] ;
   wire \mult_19_3/FS_1/C[1][2][0] ;
   wire \mult_19_3/FS_1/C[1][2][1] ;
   wire \mult_19_3/FS_1/C[1][2][2] ;
   wire \mult_19_3/FS_1/C[1][2][3] ;
   wire \mult_19_3/FS_1/C[1][3][0] ;
   wire \mult_19_3/FS_1/C[1][3][1] ;
   wire \mult_19_3/FS_1/P[0][0][1] ;
   wire \mult_19_3/FS_1/P[0][0][2] ;
   wire \mult_19_3/FS_1/P[0][0][3] ;
   wire \mult_19_3/FS_1/P[0][1][1] ;
   wire \mult_19_3/FS_1/P[0][1][2] ;
   wire \mult_19_3/FS_1/P[0][1][3] ;
   wire \mult_19_3/FS_1/P[0][2][1] ;
   wire \mult_19_3/FS_1/P[0][2][2] ;
   wire \mult_19_3/FS_1/P[0][2][3] ;
   wire \mult_19_3/FS_1/P[0][3][1] ;
   wire \mult_19_3/FS_1/TEMP_P[0][0][0] ;
   wire \mult_19_3/FS_1/TEMP_P[0][1][0] ;
   wire \mult_19_3/FS_1/TEMP_P[0][2][0] ;
   wire \mult_19_3/FS_1/TEMP_P[0][2][1] ;
   wire \mult_19_3/FS_1/TEMP_P[0][2][2] ;
   wire \mult_19_3/FS_1/TEMP_P[0][3][0] ;
   wire \mult_19_3/FS_1/G[1][0][1] ;
   wire \mult_19_3/FS_1/G[1][0][2] ;
   wire \mult_19_3/FS_1/TEMP_G[0][2][1] ;
   wire \mult_19_3/FS_1/TEMP_G[0][2][2] ;
   wire \mult_19_3/FS_1/G_n_int[0][1][3] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][0] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][1] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][2] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][3] ;
   wire \mult_19_3/FS_1/G_n_int[0][3][0] ;
   wire \mult_19_3/FS_1/PG_int[0][2][0] ;
   wire \mult_19_3/FS_1/PG_int[0][2][1] ;
   wire \mult_19_3/FS_1/PG_int[0][2][2] ;
   wire \mult_19_3/FS_1/PG_int[0][2][3] ;
   wire \mult_19_3/FS_1/PG_int[0][3][0] ;
   wire \mult_19_3/FS_1/PG_int[0][3][1] ;
   wire \mult_19_3/A2[7] ;
   wire \mult_19_3/A2[8] ;
   wire \mult_19_3/A2[9] ;
   wire \mult_19_3/A2[10] ;
   wire \mult_19_3/A2[11] ;
   wire \mult_19_3/A2[12] ;
   wire \mult_19_3/A2[13] ;
   wire \mult_19_3/A1[0] ;
   wire \mult_19_3/A1[1] ;
   wire \mult_19_3/A1[2] ;
   wire \mult_19_3/A1[3] ;
   wire \mult_19_3/A1[4] ;
   wire \mult_19_3/A1[5] ;
   wire \mult_19_3/A1[6] ;
   wire \mult_19_3/A1[7] ;
   wire \mult_19_3/A1[8] ;
   wire \mult_19_3/A1[9] ;
   wire \mult_19_3/A1[10] ;
   wire \mult_19_3/A1[11] ;
   wire \mult_19_3/A1[12] ;
   wire \mult_19_3/ab[0][1] ;
   wire \mult_19_3/ab[0][2] ;
   wire \mult_19_3/ab[0][3] ;
   wire \mult_19_3/ab[0][4] ;
   wire \mult_19_3/ab[0][5] ;
   wire \mult_19_3/ab[0][6] ;
   wire \mult_19_3/ab[0][7] ;
   wire \mult_19_3/ab[1][0] ;
   wire \mult_19_3/ab[1][1] ;
   wire \mult_19_3/ab[1][2] ;
   wire \mult_19_3/ab[1][3] ;
   wire \mult_19_3/ab[1][4] ;
   wire \mult_19_3/ab[1][5] ;
   wire \mult_19_3/ab[1][6] ;
   wire \mult_19_3/ab[1][7] ;
   wire \mult_19_3/ab[2][0] ;
   wire \mult_19_3/ab[2][1] ;
   wire \mult_19_3/ab[2][2] ;
   wire \mult_19_3/ab[2][3] ;
   wire \mult_19_3/ab[2][4] ;
   wire \mult_19_3/ab[2][5] ;
   wire \mult_19_3/ab[2][6] ;
   wire \mult_19_3/ab[2][7] ;
   wire \mult_19_3/ab[3][0] ;
   wire \mult_19_3/ab[3][1] ;
   wire \mult_19_3/ab[3][2] ;
   wire \mult_19_3/ab[3][3] ;
   wire \mult_19_3/ab[3][4] ;
   wire \mult_19_3/ab[3][5] ;
   wire \mult_19_3/ab[3][6] ;
   wire \mult_19_3/ab[3][7] ;
   wire \mult_19_3/ab[4][0] ;
   wire \mult_19_3/ab[4][1] ;
   wire \mult_19_3/ab[4][2] ;
   wire \mult_19_3/ab[4][3] ;
   wire \mult_19_3/ab[4][4] ;
   wire \mult_19_3/ab[4][5] ;
   wire \mult_19_3/ab[4][6] ;
   wire \mult_19_3/ab[4][7] ;
   wire \mult_19_3/ab[5][0] ;
   wire \mult_19_3/ab[5][1] ;
   wire \mult_19_3/ab[5][2] ;
   wire \mult_19_3/ab[5][3] ;
   wire \mult_19_3/ab[5][4] ;
   wire \mult_19_3/ab[5][5] ;
   wire \mult_19_3/ab[5][6] ;
   wire \mult_19_3/ab[5][7] ;
   wire \mult_19_3/ab[6][0] ;
   wire \mult_19_3/ab[6][1] ;
   wire \mult_19_3/ab[6][2] ;
   wire \mult_19_3/ab[6][3] ;
   wire \mult_19_3/ab[6][4] ;
   wire \mult_19_3/ab[6][5] ;
   wire \mult_19_3/ab[6][6] ;
   wire \mult_19_3/ab[6][7] ;
   wire \mult_19_3/ab[7][0] ;
   wire \mult_19_3/ab[7][1] ;
   wire \mult_19_3/ab[7][2] ;
   wire \mult_19_3/ab[7][3] ;
   wire \mult_19_3/ab[7][4] ;
   wire \mult_19_3/ab[7][5] ;
   wire \mult_19_3/ab[7][6] ;
   wire \mult_19_3/ab[7][7] ;
   wire \mult_19_3/B_not[7] ;
   wire \mult_19_3/A_not[7] ;
   wire \mult_19_2/FS_1/C[1][2][0] ;
   wire \mult_19_2/FS_1/C[1][2][1] ;
   wire \mult_19_2/FS_1/C[1][2][2] ;
   wire \mult_19_2/FS_1/C[1][2][3] ;
   wire \mult_19_2/FS_1/C[1][3][0] ;
   wire \mult_19_2/FS_1/C[1][3][1] ;
   wire \mult_19_2/FS_1/P[0][0][1] ;
   wire \mult_19_2/FS_1/P[0][0][2] ;
   wire \mult_19_2/FS_1/P[0][0][3] ;
   wire \mult_19_2/FS_1/P[0][1][1] ;
   wire \mult_19_2/FS_1/P[0][1][2] ;
   wire \mult_19_2/FS_1/P[0][1][3] ;
   wire \mult_19_2/FS_1/P[0][2][1] ;
   wire \mult_19_2/FS_1/P[0][2][2] ;
   wire \mult_19_2/FS_1/P[0][2][3] ;
   wire \mult_19_2/FS_1/P[0][3][1] ;
   wire \mult_19_2/FS_1/TEMP_P[0][0][0] ;
   wire \mult_19_2/FS_1/TEMP_P[0][1][0] ;
   wire \mult_19_2/FS_1/TEMP_P[0][2][0] ;
   wire \mult_19_2/FS_1/TEMP_P[0][2][1] ;
   wire \mult_19_2/FS_1/TEMP_P[0][2][2] ;
   wire \mult_19_2/FS_1/TEMP_P[0][3][0] ;
   wire \mult_19_2/FS_1/G[1][0][1] ;
   wire \mult_19_2/FS_1/G[1][0][2] ;
   wire \mult_19_2/FS_1/TEMP_G[0][2][1] ;
   wire \mult_19_2/FS_1/TEMP_G[0][2][2] ;
   wire \mult_19_2/FS_1/G_n_int[0][1][3] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][0] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][1] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][2] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][3] ;
   wire \mult_19_2/FS_1/G_n_int[0][3][0] ;
   wire \mult_19_2/FS_1/PG_int[0][2][0] ;
   wire \mult_19_2/FS_1/PG_int[0][2][1] ;
   wire \mult_19_2/FS_1/PG_int[0][2][2] ;
   wire \mult_19_2/FS_1/PG_int[0][2][3] ;
   wire \mult_19_2/FS_1/PG_int[0][3][0] ;
   wire \mult_19_2/FS_1/PG_int[0][3][1] ;
   wire \mult_19_2/A2[7] ;
   wire \mult_19_2/A2[8] ;
   wire \mult_19_2/A2[9] ;
   wire \mult_19_2/A2[10] ;
   wire \mult_19_2/A2[11] ;
   wire \mult_19_2/A2[12] ;
   wire \mult_19_2/A2[13] ;
   wire \mult_19_2/A1[0] ;
   wire \mult_19_2/A1[1] ;
   wire \mult_19_2/A1[2] ;
   wire \mult_19_2/A1[3] ;
   wire \mult_19_2/A1[4] ;
   wire \mult_19_2/A1[5] ;
   wire \mult_19_2/A1[6] ;
   wire \mult_19_2/A1[7] ;
   wire \mult_19_2/A1[8] ;
   wire \mult_19_2/A1[9] ;
   wire \mult_19_2/A1[10] ;
   wire \mult_19_2/A1[11] ;
   wire \mult_19_2/A1[12] ;
   wire \mult_19_2/ab[0][1] ;
   wire \mult_19_2/ab[0][2] ;
   wire \mult_19_2/ab[0][3] ;
   wire \mult_19_2/ab[0][4] ;
   wire \mult_19_2/ab[0][5] ;
   wire \mult_19_2/ab[0][6] ;
   wire \mult_19_2/ab[0][7] ;
   wire \mult_19_2/ab[1][0] ;
   wire \mult_19_2/ab[1][1] ;
   wire \mult_19_2/ab[1][2] ;
   wire \mult_19_2/ab[1][3] ;
   wire \mult_19_2/ab[1][4] ;
   wire \mult_19_2/ab[1][5] ;
   wire \mult_19_2/ab[1][6] ;
   wire \mult_19_2/ab[1][7] ;
   wire \mult_19_2/ab[2][0] ;
   wire \mult_19_2/ab[2][1] ;
   wire \mult_19_2/ab[2][2] ;
   wire \mult_19_2/ab[2][3] ;
   wire \mult_19_2/ab[2][4] ;
   wire \mult_19_2/ab[2][5] ;
   wire \mult_19_2/ab[2][6] ;
   wire \mult_19_2/ab[2][7] ;
   wire \mult_19_2/ab[3][0] ;
   wire \mult_19_2/ab[3][1] ;
   wire \mult_19_2/ab[3][2] ;
   wire \mult_19_2/ab[3][3] ;
   wire \mult_19_2/ab[3][4] ;
   wire \mult_19_2/ab[3][5] ;
   wire \mult_19_2/ab[3][6] ;
   wire \mult_19_2/ab[3][7] ;
   wire \mult_19_2/ab[4][0] ;
   wire \mult_19_2/ab[4][1] ;
   wire \mult_19_2/ab[4][2] ;
   wire \mult_19_2/ab[4][3] ;
   wire \mult_19_2/ab[4][4] ;
   wire \mult_19_2/ab[4][5] ;
   wire \mult_19_2/ab[4][6] ;
   wire \mult_19_2/ab[4][7] ;
   wire \mult_19_2/ab[5][0] ;
   wire \mult_19_2/ab[5][1] ;
   wire \mult_19_2/ab[5][2] ;
   wire \mult_19_2/ab[5][3] ;
   wire \mult_19_2/ab[5][4] ;
   wire \mult_19_2/ab[5][5] ;
   wire \mult_19_2/ab[5][6] ;
   wire \mult_19_2/ab[5][7] ;
   wire \mult_19_2/ab[6][0] ;
   wire \mult_19_2/ab[6][1] ;
   wire \mult_19_2/ab[6][2] ;
   wire \mult_19_2/ab[6][3] ;
   wire \mult_19_2/ab[6][4] ;
   wire \mult_19_2/ab[6][5] ;
   wire \mult_19_2/ab[6][6] ;
   wire \mult_19_2/ab[6][7] ;
   wire \mult_19_2/ab[7][0] ;
   wire \mult_19_2/ab[7][1] ;
   wire \mult_19_2/ab[7][2] ;
   wire \mult_19_2/ab[7][3] ;
   wire \mult_19_2/ab[7][4] ;
   wire \mult_19_2/ab[7][5] ;
   wire \mult_19_2/ab[7][6] ;
   wire \mult_19_2/ab[7][7] ;
   wire \mult_19_2/B_not[7] ;
   wire \mult_19_2/A_not[7] ;
   wire \mult_19/FS_1/C[1][2][0] ;
   wire \mult_19/FS_1/C[1][2][1] ;
   wire \mult_19/FS_1/C[1][2][2] ;
   wire \mult_19/FS_1/C[1][2][3] ;
   wire \mult_19/FS_1/C[1][3][0] ;
   wire \mult_19/FS_1/C[1][3][1] ;
   wire \mult_19/FS_1/P[0][0][1] ;
   wire \mult_19/FS_1/P[0][0][2] ;
   wire \mult_19/FS_1/P[0][0][3] ;
   wire \mult_19/FS_1/P[0][1][1] ;
   wire \mult_19/FS_1/P[0][1][2] ;
   wire \mult_19/FS_1/P[0][1][3] ;
   wire \mult_19/FS_1/P[0][2][1] ;
   wire \mult_19/FS_1/P[0][2][2] ;
   wire \mult_19/FS_1/P[0][2][3] ;
   wire \mult_19/FS_1/P[0][3][1] ;
   wire \mult_19/FS_1/TEMP_P[0][0][0] ;
   wire \mult_19/FS_1/TEMP_P[0][1][0] ;
   wire \mult_19/FS_1/TEMP_P[0][2][0] ;
   wire \mult_19/FS_1/TEMP_P[0][2][1] ;
   wire \mult_19/FS_1/TEMP_P[0][2][2] ;
   wire \mult_19/FS_1/TEMP_P[0][3][0] ;
   wire \mult_19/FS_1/G[1][0][1] ;
   wire \mult_19/FS_1/G[1][0][2] ;
   wire \mult_19/FS_1/TEMP_G[0][2][1] ;
   wire \mult_19/FS_1/TEMP_G[0][2][2] ;
   wire \mult_19/FS_1/G_n_int[0][1][3] ;
   wire \mult_19/FS_1/G_n_int[0][2][0] ;
   wire \mult_19/FS_1/G_n_int[0][2][1] ;
   wire \mult_19/FS_1/G_n_int[0][2][2] ;
   wire \mult_19/FS_1/G_n_int[0][2][3] ;
   wire \mult_19/FS_1/G_n_int[0][3][0] ;
   wire \mult_19/FS_1/PG_int[0][2][0] ;
   wire \mult_19/FS_1/PG_int[0][2][1] ;
   wire \mult_19/FS_1/PG_int[0][2][2] ;
   wire \mult_19/FS_1/PG_int[0][2][3] ;
   wire \mult_19/FS_1/PG_int[0][3][0] ;
   wire \mult_19/FS_1/PG_int[0][3][1] ;
   wire \mult_19/A2[7] ;
   wire \mult_19/A2[8] ;
   wire \mult_19/A2[9] ;
   wire \mult_19/A2[10] ;
   wire \mult_19/A2[11] ;
   wire \mult_19/A2[12] ;
   wire \mult_19/A2[13] ;
   wire \mult_19/A1[0] ;
   wire \mult_19/A1[1] ;
   wire \mult_19/A1[2] ;
   wire \mult_19/A1[3] ;
   wire \mult_19/A1[4] ;
   wire \mult_19/A1[5] ;
   wire \mult_19/A1[6] ;
   wire \mult_19/A1[7] ;
   wire \mult_19/A1[8] ;
   wire \mult_19/A1[9] ;
   wire \mult_19/A1[10] ;
   wire \mult_19/A1[11] ;
   wire \mult_19/A1[12] ;
   wire \mult_19/ab[0][1] ;
   wire \mult_19/ab[0][2] ;
   wire \mult_19/ab[0][3] ;
   wire \mult_19/ab[0][4] ;
   wire \mult_19/ab[0][5] ;
   wire \mult_19/ab[0][6] ;
   wire \mult_19/ab[0][7] ;
   wire \mult_19/ab[1][0] ;
   wire \mult_19/ab[1][1] ;
   wire \mult_19/ab[1][2] ;
   wire \mult_19/ab[1][3] ;
   wire \mult_19/ab[1][4] ;
   wire \mult_19/ab[1][5] ;
   wire \mult_19/ab[1][6] ;
   wire \mult_19/ab[1][7] ;
   wire \mult_19/ab[2][0] ;
   wire \mult_19/ab[2][1] ;
   wire \mult_19/ab[2][2] ;
   wire \mult_19/ab[2][3] ;
   wire \mult_19/ab[2][4] ;
   wire \mult_19/ab[2][5] ;
   wire \mult_19/ab[2][6] ;
   wire \mult_19/ab[2][7] ;
   wire \mult_19/ab[3][0] ;
   wire \mult_19/ab[3][1] ;
   wire \mult_19/ab[3][2] ;
   wire \mult_19/ab[3][3] ;
   wire \mult_19/ab[3][4] ;
   wire \mult_19/ab[3][5] ;
   wire \mult_19/ab[3][6] ;
   wire \mult_19/ab[3][7] ;
   wire \mult_19/ab[4][0] ;
   wire \mult_19/ab[4][1] ;
   wire \mult_19/ab[4][2] ;
   wire \mult_19/ab[4][3] ;
   wire \mult_19/ab[4][4] ;
   wire \mult_19/ab[4][5] ;
   wire \mult_19/ab[4][6] ;
   wire \mult_19/ab[4][7] ;
   wire \mult_19/ab[5][0] ;
   wire \mult_19/ab[5][1] ;
   wire \mult_19/ab[5][2] ;
   wire \mult_19/ab[5][3] ;
   wire \mult_19/ab[5][4] ;
   wire \mult_19/ab[5][5] ;
   wire \mult_19/ab[5][6] ;
   wire \mult_19/ab[5][7] ;
   wire \mult_19/ab[6][0] ;
   wire \mult_19/ab[6][1] ;
   wire \mult_19/ab[6][2] ;
   wire \mult_19/ab[6][3] ;
   wire \mult_19/ab[6][4] ;
   wire \mult_19/ab[6][5] ;
   wire \mult_19/ab[6][6] ;
   wire \mult_19/ab[6][7] ;
   wire \mult_19/ab[7][0] ;
   wire \mult_19/ab[7][1] ;
   wire \mult_19/ab[7][2] ;
   wire \mult_19/ab[7][3] ;
   wire \mult_19/ab[7][4] ;
   wire \mult_19/ab[7][5] ;
   wire \mult_19/ab[7][6] ;
   wire \mult_19/ab[7][7] ;
   wire \mult_19/B_not[7] ;
   wire \mult_19/A_not[7] ;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire [6:0] \mult_21_3/A_notx ;
   wire [6:0] \mult_21_3/B_notx ;
   wire [6:0] \mult_21_2/A_notx ;
   wire [6:0] \mult_21_2/B_notx ;
   wire [6:0] \mult_21/A_notx ;
   wire [6:0] \mult_21/B_notx ;
   wire [6:0] \mult_20_3/A_notx ;
   wire [6:0] \mult_20_3/B_notx ;
   wire [6:0] \mult_20_2/A_notx ;
   wire [6:0] \mult_20_2/B_notx ;
   wire [6:0] \mult_20/A_notx ;
   wire [6:0] \mult_20/B_notx ;
   wire [6:0] \mult_19_3/A_notx ;
   wire [6:0] \mult_19_3/B_notx ;
   wire [6:0] \mult_19_2/A_notx ;
   wire [6:0] \mult_19_2/B_notx ;
   wire [6:0] \mult_19/A_notx ;
   wire [6:0] \mult_19/B_notx ;

   inverter I_0 (.IN(rst_n),
	.OUT(N0));
   dff \result_1_reg[15]  (.D(N160),
	.CLK(n53),
	.R(N0),
	.Q(result_1[15]));
   dff \result_1_reg[14]  (.D(N159),
	.CLK(n32),
	.R(n54),
	.Q(result_1[14]));
   dff \result_1_reg[13]  (.D(N158),
	.CLK(n21),
	.R(n55),
	.Q(result_1[13]));
   dff \result_1_reg[12]  (.D(N157),
	.CLK(n39),
	.R(N0),
	.Q(result_1[12]));
   dff \result_1_reg[11]  (.D(N156),
	.CLK(n61),
	.R(n54),
	.Q(result_1[11]));
   dff \result_1_reg[10]  (.D(N155),
	.CLK(n1),
	.R(n55),
	.Q(result_1[10]));
   dff \result_1_reg[9]  (.D(N154),
	.CLK(n43),
	.R(N0),
	.Q(result_1[9]));
   dff \result_1_reg[8]  (.D(N153),
	.CLK(n47),
	.R(n54),
	.Q(result_1[8]));
   dff \result_1_reg[7]  (.D(N152),
	.CLK(n52),
	.R(n55),
	.Q(result_1[7]));
   dff \result_1_reg[6]  (.D(N151),
	.CLK(n17),
	.R(N0),
	.Q(result_1[6]));
   dff \result_1_reg[5]  (.D(N150),
	.CLK(n45),
	.R(n54),
	.Q(result_1[5]));
   dff \result_1_reg[4]  (.D(N149),
	.CLK(n44),
	.R(n55),
	.Q(result_1[4]));
   dff \result_1_reg[3]  (.D(N148),
	.CLK(n40),
	.R(N0),
	.Q(result_1[3]));
   dff \result_1_reg[2]  (.D(N147),
	.CLK(n23),
	.R(n54),
	.Q(result_1[2]));
   dff \result_1_reg[1]  (.D(N146),
	.CLK(n38),
	.R(n55),
	.Q(result_1[1]));
   dff \result_1_reg[0]  (.D(N145),
	.CLK(n34),
	.R(N0),
	.Q(result_1[0]));
   dff \result_2_reg[15]  (.D(N240),
	.CLK(n28),
	.R(n54),
	.Q(result_2[15]));
   dff \result_2_reg[14]  (.D(N239),
	.CLK(n25),
	.R(n55),
	.Q(result_2[14]));
   dff \result_2_reg[13]  (.D(N238),
	.CLK(n20),
	.R(N0),
	.Q(result_2[13]));
   dff \result_2_reg[12]  (.D(N237),
	.CLK(n22),
	.R(n54),
	.Q(result_2[12]));
   dff \result_2_reg[11]  (.D(N236),
	.CLK(n57),
	.R(n55),
	.Q(result_2[11]));
   dff \result_2_reg[10]  (.D(N235),
	.CLK(n60),
	.R(N0),
	.Q(result_2[10]));
   dff \result_2_reg[9]  (.D(N234),
	.CLK(n58),
	.R(n54),
	.Q(result_2[9]));
   dff \result_2_reg[8]  (.D(N233),
	.CLK(n29),
	.R(n55),
	.Q(result_2[8]));
   dff \result_2_reg[7]  (.D(N232),
	.CLK(n18),
	.R(N0),
	.Q(result_2[7]));
   dff \result_2_reg[6]  (.D(N231),
	.CLK(n27),
	.R(n54),
	.Q(result_2[6]));
   dff \result_2_reg[5]  (.D(N230),
	.CLK(n37),
	.R(n55),
	.Q(result_2[5]));
   dff \result_2_reg[4]  (.D(N229),
	.CLK(n65),
	.R(N0),
	.Q(result_2[4]));
   dff \result_2_reg[3]  (.D(N228),
	.CLK(n36),
	.R(n54),
	.Q(result_2[3]));
   dff \result_2_reg[2]  (.D(N227),
	.CLK(n19),
	.R(n55),
	.Q(result_2[2]));
   dff \result_2_reg[1]  (.D(N226),
	.CLK(n41),
	.R(N0),
	.Q(result_2[1]));
   dff \result_2_reg[0]  (.D(N225),
	.CLK(n26),
	.R(n54),
	.Q(result_2[0]));
   dff \result_0_reg[15]  (.D(N80),
	.CLK(n24),
	.R(n55),
	.Q(result_0[15]));
   dff \result_0_reg[14]  (.D(N79),
	.CLK(n42),
	.R(N0),
	.Q(result_0[14]));
   dff \result_0_reg[13]  (.D(N78),
	.CLK(n50),
	.R(n54),
	.Q(result_0[13]));
   dff \result_0_reg[12]  (.D(N77),
	.CLK(n63),
	.R(n55),
	.Q(result_0[12]));
   dff \result_0_reg[11]  (.D(N76),
	.CLK(n59),
	.R(N0),
	.Q(result_0[11]));
   dff \result_0_reg[10]  (.D(N75),
	.CLK(n35),
	.R(n54),
	.Q(result_0[10]));
   dff \result_0_reg[9]  (.D(N74),
	.CLK(n31),
	.R(n55),
	.Q(result_0[9]));
   dff \result_0_reg[8]  (.D(N73),
	.CLK(n30),
	.R(N0),
	.Q(result_0[8]));
   dff \result_0_reg[7]  (.D(N72),
	.CLK(n49),
	.R(n54),
	.Q(result_0[7]));
   dff \result_0_reg[6]  (.D(N71),
	.CLK(n51),
	.R(n55),
	.Q(result_0[6]));
   dff \result_0_reg[5]  (.D(N70),
	.CLK(n46),
	.R(N0),
	.Q(result_0[5]));
   dff \result_0_reg[4]  (.D(N69),
	.CLK(n64),
	.R(n54),
	.Q(result_0[4]));
   dff \result_0_reg[3]  (.D(N68),
	.CLK(n48),
	.R(n55),
	.Q(result_0[3]));
   dff \result_0_reg[2]  (.D(N67),
	.CLK(n56),
	.R(N0),
	.Q(result_0[2]));
   dff \result_0_reg[1]  (.D(N66),
	.CLK(n62),
	.R(n54),
	.Q(result_0[1]));
   dff \result_0_reg[0]  (.D(N65),
	.CLK(n33),
	.R(n55),
	.Q(result_0[0]));
   inverter U3 (.IN(clk),
	.OUT(n1));
   OAI21 \mult_21_3/FS_1/U6_1_0_3  (.OUT(\mult_21_3/FS_1/C[1][3][0] ),
	.C(n3275),
	.B(n3274),
	.A(n3273));
   OAI21 \mult_21_3/FS_1/U6_0_3_1  (.OUT(\mult_21_3/FS_1/C[1][3][1] ),
	.C(\mult_21_3/FS_1/G_n_int[0][3][0] ),
	.B(n3271),
	.A(n3270));
   XOR2 \mult_21_3/FS_1/U3_C_0_3_1  (.A(\mult_21_3/FS_1/PG_int[0][3][1] ),
	.B(\mult_21_3/FS_1/C[1][3][1] ),
	.OUT(N224));
   XOR2 \mult_21_3/FS_1/U3_C_0_3_0  (.A(\mult_21_3/FS_1/PG_int[0][3][0] ),
	.B(\mult_21_3/FS_1/C[1][3][0] ),
	.OUT(N223));
   NAND2 \mult_21_3/FS_1/U3_B_0_3_0  (.A(\mult_21_3/FS_1/G_n_int[0][3][0] ),
	.B(\mult_21_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3267));
   NAND2 \mult_21_3/FS_1/U2_0_3_0  (.A(\mult_21_3/A1[12] ),
	.B(\mult_21_3/A2[12] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_21_3/FS_1/U1_0_3_0  (.A(n3265),
	.B(n3266),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_21_3/FS_1/U6_0_2_3  (.OUT(\mult_21_3/FS_1/C[1][2][3] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][2] ),
	.B(n3264),
	.A(n3263));
   OAI21 \mult_21_3/FS_1/U5_0_2_3  (.OUT(\mult_21_3/FS_1/G[1][0][2] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][3] ),
	.B(n3262),
	.A(n3261));
   NAND2 \mult_21_3/FS_1/U4_0_2_3  (.A(\mult_21_3/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_21_3/FS_1/P[0][2][3] ),
	.OUT(n3274));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_3  (.A(\mult_21_3/FS_1/PG_int[0][2][3] ),
	.B(\mult_21_3/FS_1/C[1][2][3] ),
	.OUT(N222));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_3  (.A(\mult_21_3/FS_1/G_n_int[0][2][3] ),
	.B(\mult_21_3/FS_1/P[0][2][3] ),
	.OUT(n3260));
   NAND2 \mult_21_3/FS_1/U2_0_2_3  (.A(\mult_21_3/A1[11] ),
	.B(\mult_21_3/A2[11] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_3  (.A(n3258),
	.B(n3259),
	.OUT(\mult_21_3/FS_1/P[0][2][3] ));
   OAI21 \mult_21_3/FS_1/U6_0_2_2  (.OUT(\mult_21_3/FS_1/C[1][2][2] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][1] ),
	.B(n3257),
	.A(n3256));
   OAI21 \mult_21_3/FS_1/U5_0_2_2  (.OUT(\mult_21_3/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][2] ),
	.B(n3264),
	.A(n3255));
   NAND2 \mult_21_3/FS_1/U4_0_2_2  (.A(\mult_21_3/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_21_3/FS_1/P[0][2][2] ),
	.OUT(n3254));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_2  (.A(\mult_21_3/FS_1/PG_int[0][2][2] ),
	.B(\mult_21_3/FS_1/C[1][2][2] ),
	.OUT(N221));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_2  (.A(\mult_21_3/FS_1/G_n_int[0][2][2] ),
	.B(\mult_21_3/FS_1/P[0][2][2] ),
	.OUT(n3253));
   NAND2 \mult_21_3/FS_1/U2_0_2_2  (.A(\mult_21_3/A1[10] ),
	.B(\mult_21_3/A2[10] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_2  (.A(n3251),
	.B(n3252),
	.OUT(\mult_21_3/FS_1/P[0][2][2] ));
   OAI21 \mult_21_3/FS_1/U6_0_2_1  (.OUT(\mult_21_3/FS_1/C[1][2][1] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][0] ),
	.B(n3250),
	.A(n3273));
   OAI21 \mult_21_3/FS_1/U5_0_2_1  (.OUT(\mult_21_3/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][1] ),
	.B(n3257),
	.A(\mult_21_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_3/FS_1/U4_0_2_1  (.A(\mult_21_3/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_21_3/FS_1/P[0][2][1] ),
	.OUT(n3249));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_1  (.A(\mult_21_3/FS_1/PG_int[0][2][1] ),
	.B(\mult_21_3/FS_1/C[1][2][1] ),
	.OUT(N220));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_1  (.A(\mult_21_3/FS_1/G_n_int[0][2][1] ),
	.B(\mult_21_3/FS_1/P[0][2][1] ),
	.OUT(n3248));
   NAND2 \mult_21_3/FS_1/U2_0_2_1  (.A(\mult_21_3/A1[9] ),
	.B(\mult_21_3/A2[9] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_1  (.A(n3246),
	.B(n3247),
	.OUT(\mult_21_3/FS_1/P[0][2][1] ));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_0  (.A(\mult_21_3/FS_1/PG_int[0][2][0] ),
	.B(\mult_21_3/FS_1/C[1][2][0] ),
	.OUT(N219));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_0  (.A(\mult_21_3/FS_1/G_n_int[0][2][0] ),
	.B(\mult_21_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3245));
   NAND2 \mult_21_3/FS_1/U2_0_2_0  (.A(\mult_21_3/A1[8] ),
	.B(\mult_21_3/A2[8] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_0  (.A(n3243),
	.B(n3244),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_21_3/FS_1/U3_B_0_1_3  (.A(\mult_21_3/FS_1/G_n_int[0][1][3] ),
	.B(\mult_21_3/FS_1/P[0][1][3] ),
	.OUT(n3242));
   NAND2 \mult_21_3/FS_1/U2_0_1_3  (.A(\mult_21_3/A1[7] ),
	.B(\mult_21_3/A2[7] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_21_3/FS_1/U1_0_1_3  (.A(n3240),
	.B(n3241),
	.OUT(\mult_21_3/FS_1/P[0][1][3] ));
   inverter \mult_21_3/AN1_7  (.IN(matrix22[7]),
	.OUT(\mult_21_3/A_not[7] ));
   inverter \mult_21_3/AN1_6  (.IN(matrix22[6]),
	.OUT(\mult_21_3/A_notx [6]));
   inverter \mult_21_3/AN1_5  (.IN(matrix22[5]),
	.OUT(\mult_21_3/A_notx [5]));
   inverter \mult_21_3/AN1_4  (.IN(matrix22[4]),
	.OUT(\mult_21_3/A_notx [4]));
   inverter \mult_21_3/AN1_3  (.IN(matrix22[3]),
	.OUT(\mult_21_3/A_notx [3]));
   inverter \mult_21_3/AN1_2  (.IN(matrix22[2]),
	.OUT(\mult_21_3/A_notx [2]));
   inverter \mult_21_3/AN1_1  (.IN(matrix22[1]),
	.OUT(\mult_21_3/A_notx [1]));
   inverter \mult_21_3/AN1_0  (.IN(matrix22[0]),
	.OUT(\mult_21_3/A_notx [0]));
   inverter \mult_21_3/AN1_7_0  (.IN(vector_2[7]),
	.OUT(\mult_21_3/B_not[7] ));
   inverter \mult_21_3/AN1_6_0  (.IN(vector_2[6]),
	.OUT(\mult_21_3/B_notx [6]));
   inverter \mult_21_3/AN1_5_0  (.IN(vector_2[5]),
	.OUT(\mult_21_3/B_notx [5]));
   inverter \mult_21_3/AN1_4_0  (.IN(vector_2[4]),
	.OUT(\mult_21_3/B_notx [4]));
   inverter \mult_21_3/AN1_3_0  (.IN(vector_2[3]),
	.OUT(\mult_21_3/B_notx [3]));
   inverter \mult_21_3/AN1_2_0  (.IN(vector_2[2]),
	.OUT(\mult_21_3/B_notx [2]));
   inverter \mult_21_3/AN1_1_0  (.IN(vector_2[1]),
	.OUT(\mult_21_3/B_notx [1]));
   inverter \mult_21_3/AN1_0_0  (.IN(vector_2[0]),
	.OUT(\mult_21_3/B_notx [0]));
   NOR2 \mult_21_3/AN1_7_7  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[7][7] ));
   NOR2 \mult_21_3/AN3_7_6  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[7][6] ));
   NOR2 \mult_21_3/AN3_7_5  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[7][5] ));
   NOR2 \mult_21_3/AN3_7_4  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[7][4] ));
   NOR2 \mult_21_3/AN3_7_3  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[7][3] ));
   NOR2 \mult_21_3/AN3_7_2  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[7][2] ));
   NOR2 \mult_21_3/AN3_7_1  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[7][1] ));
   NOR2 \mult_21_3/AN3_7_0  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[7][0] ));
   NOR2 \mult_21_3/AN2_6_7  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[6][7] ));
   NOR2 \mult_21_3/AN1_6_6  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[6][6] ));
   NOR2 \mult_21_3/AN1_6_5  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[6][5] ));
   NOR2 \mult_21_3/AN1_6_4  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[6][4] ));
   NOR2 \mult_21_3/AN1_6_3  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[6][3] ));
   NOR2 \mult_21_3/AN1_6_2  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[6][2] ));
   NOR2 \mult_21_3/AN1_6_1  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[6][1] ));
   NOR2 \mult_21_3/AN1_6_0_0  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[6][0] ));
   NOR2 \mult_21_3/AN2_5_7  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[5][7] ));
   NOR2 \mult_21_3/AN1_5_6  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[5][6] ));
   NOR2 \mult_21_3/AN1_5_5  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[5][5] ));
   NOR2 \mult_21_3/AN1_5_4  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[5][4] ));
   NOR2 \mult_21_3/AN1_5_3  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[5][3] ));
   NOR2 \mult_21_3/AN1_5_2  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[5][2] ));
   NOR2 \mult_21_3/AN1_5_1  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[5][1] ));
   NOR2 \mult_21_3/AN1_5_0_0  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[5][0] ));
   NOR2 \mult_21_3/AN2_4_7  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[4][7] ));
   NOR2 \mult_21_3/AN1_4_6  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[4][6] ));
   NOR2 \mult_21_3/AN1_4_5  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[4][5] ));
   NOR2 \mult_21_3/AN1_4_4  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[4][4] ));
   NOR2 \mult_21_3/AN1_4_3  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[4][3] ));
   NOR2 \mult_21_3/AN1_4_2  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[4][2] ));
   NOR2 \mult_21_3/AN1_4_1  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[4][1] ));
   NOR2 \mult_21_3/AN1_4_0_0  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[4][0] ));
   NOR2 \mult_21_3/AN2_3_7  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[3][7] ));
   NOR2 \mult_21_3/AN1_3_6  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[3][6] ));
   NOR2 \mult_21_3/AN1_3_5  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[3][5] ));
   NOR2 \mult_21_3/AN1_3_4  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[3][4] ));
   NOR2 \mult_21_3/AN1_3_3  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[3][3] ));
   NOR2 \mult_21_3/AN1_3_2  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[3][2] ));
   NOR2 \mult_21_3/AN1_3_1  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[3][1] ));
   NOR2 \mult_21_3/AN1_3_0_0  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[3][0] ));
   NOR2 \mult_21_3/AN2_2_7  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[2][7] ));
   NOR2 \mult_21_3/AN1_2_6  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[2][6] ));
   NOR2 \mult_21_3/AN1_2_5  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[2][5] ));
   NOR2 \mult_21_3/AN1_2_4  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[2][4] ));
   NOR2 \mult_21_3/AN1_2_3  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[2][3] ));
   NOR2 \mult_21_3/AN1_2_2  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[2][2] ));
   NOR2 \mult_21_3/AN1_2_1  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[2][1] ));
   NOR2 \mult_21_3/AN1_2_0_0  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[2][0] ));
   NOR2 \mult_21_3/AN2_1_7  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[1][7] ));
   NOR2 \mult_21_3/AN1_1_6  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[1][6] ));
   NOR2 \mult_21_3/AN1_1_5  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[1][5] ));
   NOR2 \mult_21_3/AN1_1_4  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[1][4] ));
   NOR2 \mult_21_3/AN1_1_3  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[1][3] ));
   NOR2 \mult_21_3/AN1_1_2  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[1][2] ));
   NOR2 \mult_21_3/AN1_1_1  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[1][1] ));
   NOR2 \mult_21_3/AN1_1_0_0  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[1][0] ));
   NOR2 \mult_21_3/AN2_0_7  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[0][7] ));
   NOR2 \mult_21_3/AN1_0_6  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[0][6] ));
   NOR2 \mult_21_3/AN1_0_5  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[0][5] ));
   NOR2 \mult_21_3/AN1_0_4  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[0][4] ));
   NOR2 \mult_21_3/AN1_0_3  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[0][3] ));
   NOR2 \mult_21_3/AN1_0_2  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[0][2] ));
   NOR2 \mult_21_3/AN1_0_1  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[0][1] ));
   NOR2 \mult_21_3/AN1_0_0_0  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(N209));
   OAI21 \mult_21_2/FS_1/U6_1_0_3  (.OUT(\mult_21_2/FS_1/C[1][3][0] ),
	.C(n3225),
	.B(n3224),
	.A(n3223));
   OAI21 \mult_21_2/FS_1/U6_0_3_1  (.OUT(\mult_21_2/FS_1/C[1][3][1] ),
	.C(\mult_21_2/FS_1/G_n_int[0][3][0] ),
	.B(n3221),
	.A(n3220));
   XOR2 \mult_21_2/FS_1/U3_C_0_3_1  (.A(\mult_21_2/FS_1/PG_int[0][3][1] ),
	.B(\mult_21_2/FS_1/C[1][3][1] ),
	.OUT(N192));
   XOR2 \mult_21_2/FS_1/U3_C_0_3_0  (.A(\mult_21_2/FS_1/PG_int[0][3][0] ),
	.B(\mult_21_2/FS_1/C[1][3][0] ),
	.OUT(N191));
   NAND2 \mult_21_2/FS_1/U3_B_0_3_0  (.A(\mult_21_2/FS_1/G_n_int[0][3][0] ),
	.B(\mult_21_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3217));
   NAND2 \mult_21_2/FS_1/U2_0_3_0  (.A(\mult_21_2/A1[12] ),
	.B(\mult_21_2/A2[12] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_21_2/FS_1/U1_0_3_0  (.A(n3215),
	.B(n3216),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_21_2/FS_1/U6_0_2_3  (.OUT(\mult_21_2/FS_1/C[1][2][3] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][2] ),
	.B(n3214),
	.A(n3213));
   OAI21 \mult_21_2/FS_1/U5_0_2_3  (.OUT(\mult_21_2/FS_1/G[1][0][2] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][3] ),
	.B(n3212),
	.A(n3211));
   NAND2 \mult_21_2/FS_1/U4_0_2_3  (.A(\mult_21_2/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_21_2/FS_1/P[0][2][3] ),
	.OUT(n3224));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_3  (.A(\mult_21_2/FS_1/PG_int[0][2][3] ),
	.B(\mult_21_2/FS_1/C[1][2][3] ),
	.OUT(N190));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_3  (.A(\mult_21_2/FS_1/G_n_int[0][2][3] ),
	.B(\mult_21_2/FS_1/P[0][2][3] ),
	.OUT(n3210));
   NAND2 \mult_21_2/FS_1/U2_0_2_3  (.A(\mult_21_2/A1[11] ),
	.B(\mult_21_2/A2[11] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_3  (.A(n3208),
	.B(n3209),
	.OUT(\mult_21_2/FS_1/P[0][2][3] ));
   OAI21 \mult_21_2/FS_1/U6_0_2_2  (.OUT(\mult_21_2/FS_1/C[1][2][2] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][1] ),
	.B(n3207),
	.A(n3206));
   OAI21 \mult_21_2/FS_1/U5_0_2_2  (.OUT(\mult_21_2/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][2] ),
	.B(n3214),
	.A(n3205));
   NAND2 \mult_21_2/FS_1/U4_0_2_2  (.A(\mult_21_2/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_21_2/FS_1/P[0][2][2] ),
	.OUT(n3204));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_2  (.A(\mult_21_2/FS_1/PG_int[0][2][2] ),
	.B(\mult_21_2/FS_1/C[1][2][2] ),
	.OUT(N189));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_2  (.A(\mult_21_2/FS_1/G_n_int[0][2][2] ),
	.B(\mult_21_2/FS_1/P[0][2][2] ),
	.OUT(n3203));
   NAND2 \mult_21_2/FS_1/U2_0_2_2  (.A(\mult_21_2/A1[10] ),
	.B(\mult_21_2/A2[10] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_2  (.A(n3201),
	.B(n3202),
	.OUT(\mult_21_2/FS_1/P[0][2][2] ));
   OAI21 \mult_21_2/FS_1/U6_0_2_1  (.OUT(\mult_21_2/FS_1/C[1][2][1] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][0] ),
	.B(n3200),
	.A(n3223));
   OAI21 \mult_21_2/FS_1/U5_0_2_1  (.OUT(\mult_21_2/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][1] ),
	.B(n3207),
	.A(\mult_21_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_2/FS_1/U4_0_2_1  (.A(\mult_21_2/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_21_2/FS_1/P[0][2][1] ),
	.OUT(n3199));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_1  (.A(\mult_21_2/FS_1/PG_int[0][2][1] ),
	.B(\mult_21_2/FS_1/C[1][2][1] ),
	.OUT(N188));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_1  (.A(\mult_21_2/FS_1/G_n_int[0][2][1] ),
	.B(\mult_21_2/FS_1/P[0][2][1] ),
	.OUT(n3198));
   NAND2 \mult_21_2/FS_1/U2_0_2_1  (.A(\mult_21_2/A1[9] ),
	.B(\mult_21_2/A2[9] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_1  (.A(n3196),
	.B(n3197),
	.OUT(\mult_21_2/FS_1/P[0][2][1] ));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_0  (.A(\mult_21_2/FS_1/PG_int[0][2][0] ),
	.B(\mult_21_2/FS_1/C[1][2][0] ),
	.OUT(N187));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_0  (.A(\mult_21_2/FS_1/G_n_int[0][2][0] ),
	.B(\mult_21_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3195));
   NAND2 \mult_21_2/FS_1/U2_0_2_0  (.A(\mult_21_2/A1[8] ),
	.B(\mult_21_2/A2[8] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_0  (.A(n3193),
	.B(n3194),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_21_2/FS_1/U3_B_0_1_3  (.A(\mult_21_2/FS_1/G_n_int[0][1][3] ),
	.B(\mult_21_2/FS_1/P[0][1][3] ),
	.OUT(n3192));
   NAND2 \mult_21_2/FS_1/U2_0_1_3  (.A(\mult_21_2/A1[7] ),
	.B(\mult_21_2/A2[7] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_21_2/FS_1/U1_0_1_3  (.A(n3190),
	.B(n3191),
	.OUT(\mult_21_2/FS_1/P[0][1][3] ));
   inverter \mult_21_2/AN1_7  (.IN(matrix21[7]),
	.OUT(\mult_21_2/A_not[7] ));
   inverter \mult_21_2/AN1_6  (.IN(matrix21[6]),
	.OUT(\mult_21_2/A_notx [6]));
   inverter \mult_21_2/AN1_5  (.IN(matrix21[5]),
	.OUT(\mult_21_2/A_notx [5]));
   inverter \mult_21_2/AN1_4  (.IN(matrix21[4]),
	.OUT(\mult_21_2/A_notx [4]));
   inverter \mult_21_2/AN1_3  (.IN(matrix21[3]),
	.OUT(\mult_21_2/A_notx [3]));
   inverter \mult_21_2/AN1_2  (.IN(matrix21[2]),
	.OUT(\mult_21_2/A_notx [2]));
   inverter \mult_21_2/AN1_1  (.IN(matrix21[1]),
	.OUT(\mult_21_2/A_notx [1]));
   inverter \mult_21_2/AN1_0  (.IN(matrix21[0]),
	.OUT(\mult_21_2/A_notx [0]));
   inverter \mult_21_2/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_21_2/B_not[7] ));
   inverter \mult_21_2/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_21_2/B_notx [6]));
   inverter \mult_21_2/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_21_2/B_notx [5]));
   inverter \mult_21_2/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_21_2/B_notx [4]));
   inverter \mult_21_2/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_21_2/B_notx [3]));
   inverter \mult_21_2/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_21_2/B_notx [2]));
   inverter \mult_21_2/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_21_2/B_notx [1]));
   inverter \mult_21_2/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_21_2/B_notx [0]));
   NOR2 \mult_21_2/AN1_7_7  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[7][7] ));
   NOR2 \mult_21_2/AN3_7_6  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[7][6] ));
   NOR2 \mult_21_2/AN3_7_5  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[7][5] ));
   NOR2 \mult_21_2/AN3_7_4  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[7][4] ));
   NOR2 \mult_21_2/AN3_7_3  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[7][3] ));
   NOR2 \mult_21_2/AN3_7_2  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[7][2] ));
   NOR2 \mult_21_2/AN3_7_1  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[7][1] ));
   NOR2 \mult_21_2/AN3_7_0  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[7][0] ));
   NOR2 \mult_21_2/AN2_6_7  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[6][7] ));
   NOR2 \mult_21_2/AN1_6_6  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[6][6] ));
   NOR2 \mult_21_2/AN1_6_5  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[6][5] ));
   NOR2 \mult_21_2/AN1_6_4  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[6][4] ));
   NOR2 \mult_21_2/AN1_6_3  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[6][3] ));
   NOR2 \mult_21_2/AN1_6_2  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[6][2] ));
   NOR2 \mult_21_2/AN1_6_1  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[6][1] ));
   NOR2 \mult_21_2/AN1_6_0_0  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[6][0] ));
   NOR2 \mult_21_2/AN2_5_7  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[5][7] ));
   NOR2 \mult_21_2/AN1_5_6  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[5][6] ));
   NOR2 \mult_21_2/AN1_5_5  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[5][5] ));
   NOR2 \mult_21_2/AN1_5_4  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[5][4] ));
   NOR2 \mult_21_2/AN1_5_3  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[5][3] ));
   NOR2 \mult_21_2/AN1_5_2  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[5][2] ));
   NOR2 \mult_21_2/AN1_5_1  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[5][1] ));
   NOR2 \mult_21_2/AN1_5_0_0  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[5][0] ));
   NOR2 \mult_21_2/AN2_4_7  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[4][7] ));
   NOR2 \mult_21_2/AN1_4_6  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[4][6] ));
   NOR2 \mult_21_2/AN1_4_5  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[4][5] ));
   NOR2 \mult_21_2/AN1_4_4  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[4][4] ));
   NOR2 \mult_21_2/AN1_4_3  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[4][3] ));
   NOR2 \mult_21_2/AN1_4_2  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[4][2] ));
   NOR2 \mult_21_2/AN1_4_1  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[4][1] ));
   NOR2 \mult_21_2/AN1_4_0_0  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[4][0] ));
   NOR2 \mult_21_2/AN2_3_7  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[3][7] ));
   NOR2 \mult_21_2/AN1_3_6  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[3][6] ));
   NOR2 \mult_21_2/AN1_3_5  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[3][5] ));
   NOR2 \mult_21_2/AN1_3_4  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[3][4] ));
   NOR2 \mult_21_2/AN1_3_3  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[3][3] ));
   NOR2 \mult_21_2/AN1_3_2  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[3][2] ));
   NOR2 \mult_21_2/AN1_3_1  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[3][1] ));
   NOR2 \mult_21_2/AN1_3_0_0  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[3][0] ));
   NOR2 \mult_21_2/AN2_2_7  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[2][7] ));
   NOR2 \mult_21_2/AN1_2_6  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[2][6] ));
   NOR2 \mult_21_2/AN1_2_5  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[2][5] ));
   NOR2 \mult_21_2/AN1_2_4  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[2][4] ));
   NOR2 \mult_21_2/AN1_2_3  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[2][3] ));
   NOR2 \mult_21_2/AN1_2_2  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[2][2] ));
   NOR2 \mult_21_2/AN1_2_1  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[2][1] ));
   NOR2 \mult_21_2/AN1_2_0_0  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[2][0] ));
   NOR2 \mult_21_2/AN2_1_7  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[1][7] ));
   NOR2 \mult_21_2/AN1_1_6  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[1][6] ));
   NOR2 \mult_21_2/AN1_1_5  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[1][5] ));
   NOR2 \mult_21_2/AN1_1_4  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[1][4] ));
   NOR2 \mult_21_2/AN1_1_3  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[1][3] ));
   NOR2 \mult_21_2/AN1_1_2  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[1][2] ));
   NOR2 \mult_21_2/AN1_1_1  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[1][1] ));
   NOR2 \mult_21_2/AN1_1_0_0  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[1][0] ));
   NOR2 \mult_21_2/AN2_0_7  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[0][7] ));
   NOR2 \mult_21_2/AN1_0_6  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[0][6] ));
   NOR2 \mult_21_2/AN1_0_5  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[0][5] ));
   NOR2 \mult_21_2/AN1_0_4  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[0][4] ));
   NOR2 \mult_21_2/AN1_0_3  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[0][3] ));
   NOR2 \mult_21_2/AN1_0_2  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[0][2] ));
   NOR2 \mult_21_2/AN1_0_1  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[0][1] ));
   NOR2 \mult_21_2/AN1_0_0_0  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(N177));
   OAI21 \mult_21/FS_1/U6_1_0_3  (.OUT(\mult_21/FS_1/C[1][3][0] ),
	.C(n3175),
	.B(n3174),
	.A(n3173));
   OAI21 \mult_21/FS_1/U6_0_3_1  (.OUT(\mult_21/FS_1/C[1][3][1] ),
	.C(\mult_21/FS_1/G_n_int[0][3][0] ),
	.B(n3171),
	.A(n3170));
   XOR2 \mult_21/FS_1/U3_C_0_3_1  (.A(\mult_21/FS_1/PG_int[0][3][1] ),
	.B(\mult_21/FS_1/C[1][3][1] ),
	.OUT(N176));
   XOR2 \mult_21/FS_1/U3_C_0_3_0  (.A(\mult_21/FS_1/PG_int[0][3][0] ),
	.B(\mult_21/FS_1/C[1][3][0] ),
	.OUT(N175));
   NAND2 \mult_21/FS_1/U3_B_0_3_0  (.A(\mult_21/FS_1/G_n_int[0][3][0] ),
	.B(\mult_21/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3167));
   NAND2 \mult_21/FS_1/U2_0_3_0  (.A(\mult_21/A1[12] ),
	.B(\mult_21/A2[12] ),
	.OUT(\mult_21/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_21/FS_1/U1_0_3_0  (.A(n3165),
	.B(n3166),
	.OUT(\mult_21/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_21/FS_1/U6_0_2_3  (.OUT(\mult_21/FS_1/C[1][2][3] ),
	.C(\mult_21/FS_1/G_n_int[0][2][2] ),
	.B(n3164),
	.A(n3163));
   OAI21 \mult_21/FS_1/U5_0_2_3  (.OUT(\mult_21/FS_1/G[1][0][2] ),
	.C(\mult_21/FS_1/G_n_int[0][2][3] ),
	.B(n3162),
	.A(n3161));
   NAND2 \mult_21/FS_1/U4_0_2_3  (.A(\mult_21/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_21/FS_1/P[0][2][3] ),
	.OUT(n3174));
   XOR2 \mult_21/FS_1/U3_C_0_2_3  (.A(\mult_21/FS_1/PG_int[0][2][3] ),
	.B(\mult_21/FS_1/C[1][2][3] ),
	.OUT(N174));
   NAND2 \mult_21/FS_1/U3_B_0_2_3  (.A(\mult_21/FS_1/G_n_int[0][2][3] ),
	.B(\mult_21/FS_1/P[0][2][3] ),
	.OUT(n3160));
   NAND2 \mult_21/FS_1/U2_0_2_3  (.A(\mult_21/A1[11] ),
	.B(\mult_21/A2[11] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_21/FS_1/U1_0_2_3  (.A(n3158),
	.B(n3159),
	.OUT(\mult_21/FS_1/P[0][2][3] ));
   OAI21 \mult_21/FS_1/U6_0_2_2  (.OUT(\mult_21/FS_1/C[1][2][2] ),
	.C(\mult_21/FS_1/G_n_int[0][2][1] ),
	.B(n3157),
	.A(n3156));
   OAI21 \mult_21/FS_1/U5_0_2_2  (.OUT(\mult_21/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_21/FS_1/G_n_int[0][2][2] ),
	.B(n3164),
	.A(n3155));
   NAND2 \mult_21/FS_1/U4_0_2_2  (.A(\mult_21/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_21/FS_1/P[0][2][2] ),
	.OUT(n3154));
   XOR2 \mult_21/FS_1/U3_C_0_2_2  (.A(\mult_21/FS_1/PG_int[0][2][2] ),
	.B(\mult_21/FS_1/C[1][2][2] ),
	.OUT(N173));
   NAND2 \mult_21/FS_1/U3_B_0_2_2  (.A(\mult_21/FS_1/G_n_int[0][2][2] ),
	.B(\mult_21/FS_1/P[0][2][2] ),
	.OUT(n3153));
   NAND2 \mult_21/FS_1/U2_0_2_2  (.A(\mult_21/A1[10] ),
	.B(\mult_21/A2[10] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_21/FS_1/U1_0_2_2  (.A(n3151),
	.B(n3152),
	.OUT(\mult_21/FS_1/P[0][2][2] ));
   OAI21 \mult_21/FS_1/U6_0_2_1  (.OUT(\mult_21/FS_1/C[1][2][1] ),
	.C(\mult_21/FS_1/G_n_int[0][2][0] ),
	.B(n3150),
	.A(n3173));
   OAI21 \mult_21/FS_1/U5_0_2_1  (.OUT(\mult_21/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_21/FS_1/G_n_int[0][2][1] ),
	.B(n3157),
	.A(\mult_21/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21/FS_1/U4_0_2_1  (.A(\mult_21/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_21/FS_1/P[0][2][1] ),
	.OUT(n3149));
   XOR2 \mult_21/FS_1/U3_C_0_2_1  (.A(\mult_21/FS_1/PG_int[0][2][1] ),
	.B(\mult_21/FS_1/C[1][2][1] ),
	.OUT(N172));
   NAND2 \mult_21/FS_1/U3_B_0_2_1  (.A(\mult_21/FS_1/G_n_int[0][2][1] ),
	.B(\mult_21/FS_1/P[0][2][1] ),
	.OUT(n3148));
   NAND2 \mult_21/FS_1/U2_0_2_1  (.A(\mult_21/A1[9] ),
	.B(\mult_21/A2[9] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_21/FS_1/U1_0_2_1  (.A(n3146),
	.B(n3147),
	.OUT(\mult_21/FS_1/P[0][2][1] ));
   XOR2 \mult_21/FS_1/U3_C_0_2_0  (.A(\mult_21/FS_1/PG_int[0][2][0] ),
	.B(\mult_21/FS_1/C[1][2][0] ),
	.OUT(N171));
   NAND2 \mult_21/FS_1/U3_B_0_2_0  (.A(\mult_21/FS_1/G_n_int[0][2][0] ),
	.B(\mult_21/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3145));
   NAND2 \mult_21/FS_1/U2_0_2_0  (.A(\mult_21/A1[8] ),
	.B(\mult_21/A2[8] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21/FS_1/U1_0_2_0  (.A(n3143),
	.B(n3144),
	.OUT(\mult_21/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_21/FS_1/U3_B_0_1_3  (.A(\mult_21/FS_1/G_n_int[0][1][3] ),
	.B(\mult_21/FS_1/P[0][1][3] ),
	.OUT(n3142));
   NAND2 \mult_21/FS_1/U2_0_1_3  (.A(\mult_21/A1[7] ),
	.B(\mult_21/A2[7] ),
	.OUT(\mult_21/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_21/FS_1/U1_0_1_3  (.A(n3140),
	.B(n3141),
	.OUT(\mult_21/FS_1/P[0][1][3] ));
   inverter \mult_21/AN1_7  (.IN(matrix20[7]),
	.OUT(\mult_21/A_not[7] ));
   inverter \mult_21/AN1_6  (.IN(matrix20[6]),
	.OUT(\mult_21/A_notx [6]));
   inverter \mult_21/AN1_5  (.IN(matrix20[5]),
	.OUT(\mult_21/A_notx [5]));
   inverter \mult_21/AN1_4  (.IN(matrix20[4]),
	.OUT(\mult_21/A_notx [4]));
   inverter \mult_21/AN1_3  (.IN(matrix20[3]),
	.OUT(\mult_21/A_notx [3]));
   inverter \mult_21/AN1_2  (.IN(matrix20[2]),
	.OUT(\mult_21/A_notx [2]));
   inverter \mult_21/AN1_1  (.IN(matrix20[1]),
	.OUT(\mult_21/A_notx [1]));
   inverter \mult_21/AN1_0  (.IN(matrix20[0]),
	.OUT(\mult_21/A_notx [0]));
   inverter \mult_21/AN1_7_0  (.IN(vector_0[7]),
	.OUT(\mult_21/B_not[7] ));
   inverter \mult_21/AN1_6_0  (.IN(vector_0[6]),
	.OUT(\mult_21/B_notx [6]));
   inverter \mult_21/AN1_5_0  (.IN(vector_0[5]),
	.OUT(\mult_21/B_notx [5]));
   inverter \mult_21/AN1_4_0  (.IN(vector_0[4]),
	.OUT(\mult_21/B_notx [4]));
   inverter \mult_21/AN1_3_0  (.IN(vector_0[3]),
	.OUT(\mult_21/B_notx [3]));
   inverter \mult_21/AN1_2_0  (.IN(vector_0[2]),
	.OUT(\mult_21/B_notx [2]));
   inverter \mult_21/AN1_1_0  (.IN(vector_0[1]),
	.OUT(\mult_21/B_notx [1]));
   inverter \mult_21/AN1_0_0  (.IN(vector_0[0]),
	.OUT(\mult_21/B_notx [0]));
   NOR2 \mult_21/AN1_7_7  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[7][7] ));
   NOR2 \mult_21/AN3_7_6  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[7][6] ));
   NOR2 \mult_21/AN3_7_5  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[7][5] ));
   NOR2 \mult_21/AN3_7_4  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[7][4] ));
   NOR2 \mult_21/AN3_7_3  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[7][3] ));
   NOR2 \mult_21/AN3_7_2  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[7][2] ));
   NOR2 \mult_21/AN3_7_1  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[7][1] ));
   NOR2 \mult_21/AN3_7_0  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[7][0] ));
   NOR2 \mult_21/AN2_6_7  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[6][7] ));
   NOR2 \mult_21/AN1_6_6  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[6][6] ));
   NOR2 \mult_21/AN1_6_5  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[6][5] ));
   NOR2 \mult_21/AN1_6_4  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[6][4] ));
   NOR2 \mult_21/AN1_6_3  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[6][3] ));
   NOR2 \mult_21/AN1_6_2  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[6][2] ));
   NOR2 \mult_21/AN1_6_1  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[6][1] ));
   NOR2 \mult_21/AN1_6_0_0  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[6][0] ));
   NOR2 \mult_21/AN2_5_7  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[5][7] ));
   NOR2 \mult_21/AN1_5_6  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[5][6] ));
   NOR2 \mult_21/AN1_5_5  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[5][5] ));
   NOR2 \mult_21/AN1_5_4  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[5][4] ));
   NOR2 \mult_21/AN1_5_3  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[5][3] ));
   NOR2 \mult_21/AN1_5_2  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[5][2] ));
   NOR2 \mult_21/AN1_5_1  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[5][1] ));
   NOR2 \mult_21/AN1_5_0_0  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[5][0] ));
   NOR2 \mult_21/AN2_4_7  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[4][7] ));
   NOR2 \mult_21/AN1_4_6  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[4][6] ));
   NOR2 \mult_21/AN1_4_5  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[4][5] ));
   NOR2 \mult_21/AN1_4_4  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[4][4] ));
   NOR2 \mult_21/AN1_4_3  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[4][3] ));
   NOR2 \mult_21/AN1_4_2  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[4][2] ));
   NOR2 \mult_21/AN1_4_1  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[4][1] ));
   NOR2 \mult_21/AN1_4_0_0  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[4][0] ));
   NOR2 \mult_21/AN2_3_7  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[3][7] ));
   NOR2 \mult_21/AN1_3_6  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[3][6] ));
   NOR2 \mult_21/AN1_3_5  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[3][5] ));
   NOR2 \mult_21/AN1_3_4  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[3][4] ));
   NOR2 \mult_21/AN1_3_3  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[3][3] ));
   NOR2 \mult_21/AN1_3_2  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[3][2] ));
   NOR2 \mult_21/AN1_3_1  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[3][1] ));
   NOR2 \mult_21/AN1_3_0_0  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[3][0] ));
   NOR2 \mult_21/AN2_2_7  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[2][7] ));
   NOR2 \mult_21/AN1_2_6  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[2][6] ));
   NOR2 \mult_21/AN1_2_5  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[2][5] ));
   NOR2 \mult_21/AN1_2_4  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[2][4] ));
   NOR2 \mult_21/AN1_2_3  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[2][3] ));
   NOR2 \mult_21/AN1_2_2  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[2][2] ));
   NOR2 \mult_21/AN1_2_1  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[2][1] ));
   NOR2 \mult_21/AN1_2_0_0  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[2][0] ));
   NOR2 \mult_21/AN2_1_7  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[1][7] ));
   NOR2 \mult_21/AN1_1_6  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[1][6] ));
   NOR2 \mult_21/AN1_1_5  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[1][5] ));
   NOR2 \mult_21/AN1_1_4  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[1][4] ));
   NOR2 \mult_21/AN1_1_3  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[1][3] ));
   NOR2 \mult_21/AN1_1_2  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[1][2] ));
   NOR2 \mult_21/AN1_1_1  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[1][1] ));
   NOR2 \mult_21/AN1_1_0_0  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[1][0] ));
   NOR2 \mult_21/AN2_0_7  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[0][7] ));
   NOR2 \mult_21/AN1_0_6  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[0][6] ));
   NOR2 \mult_21/AN1_0_5  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[0][5] ));
   NOR2 \mult_21/AN1_0_4  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[0][4] ));
   NOR2 \mult_21/AN1_0_3  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[0][3] ));
   NOR2 \mult_21/AN1_0_2  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[0][2] ));
   NOR2 \mult_21/AN1_0_1  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[0][1] ));
   NOR2 \mult_21/AN1_0_0_0  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [0]),
	.OUT(N161));
   OAI21 \mult_20_3/FS_1/U6_1_0_3  (.OUT(\mult_20_3/FS_1/C[1][3][0] ),
	.C(n3125),
	.B(n3124),
	.A(n3123));
   OAI21 \mult_20_3/FS_1/U6_0_3_1  (.OUT(\mult_20_3/FS_1/C[1][3][1] ),
	.C(\mult_20_3/FS_1/G_n_int[0][3][0] ),
	.B(n3121),
	.A(n3120));
   XOR2 \mult_20_3/FS_1/U3_C_0_3_1  (.A(\mult_20_3/FS_1/PG_int[0][3][1] ),
	.B(\mult_20_3/FS_1/C[1][3][1] ),
	.OUT(N144));
   XOR2 \mult_20_3/FS_1/U3_C_0_3_0  (.A(\mult_20_3/FS_1/PG_int[0][3][0] ),
	.B(\mult_20_3/FS_1/C[1][3][0] ),
	.OUT(N143));
   NAND2 \mult_20_3/FS_1/U3_B_0_3_0  (.A(\mult_20_3/FS_1/G_n_int[0][3][0] ),
	.B(\mult_20_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3117));
   NAND2 \mult_20_3/FS_1/U2_0_3_0  (.A(\mult_20_3/A1[12] ),
	.B(\mult_20_3/A2[12] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_20_3/FS_1/U1_0_3_0  (.A(n3115),
	.B(n3116),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_20_3/FS_1/U6_0_2_3  (.OUT(\mult_20_3/FS_1/C[1][2][3] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][2] ),
	.B(n3114),
	.A(n3113));
   OAI21 \mult_20_3/FS_1/U5_0_2_3  (.OUT(\mult_20_3/FS_1/G[1][0][2] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][3] ),
	.B(n3112),
	.A(n3111));
   NAND2 \mult_20_3/FS_1/U4_0_2_3  (.A(\mult_20_3/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_20_3/FS_1/P[0][2][3] ),
	.OUT(n3124));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_3  (.A(\mult_20_3/FS_1/PG_int[0][2][3] ),
	.B(\mult_20_3/FS_1/C[1][2][3] ),
	.OUT(N142));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_3  (.A(\mult_20_3/FS_1/G_n_int[0][2][3] ),
	.B(\mult_20_3/FS_1/P[0][2][3] ),
	.OUT(n3110));
   NAND2 \mult_20_3/FS_1/U2_0_2_3  (.A(\mult_20_3/A1[11] ),
	.B(\mult_20_3/A2[11] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_3  (.A(n3108),
	.B(n3109),
	.OUT(\mult_20_3/FS_1/P[0][2][3] ));
   OAI21 \mult_20_3/FS_1/U6_0_2_2  (.OUT(\mult_20_3/FS_1/C[1][2][2] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][1] ),
	.B(n3107),
	.A(n3106));
   OAI21 \mult_20_3/FS_1/U5_0_2_2  (.OUT(\mult_20_3/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][2] ),
	.B(n3114),
	.A(n3105));
   NAND2 \mult_20_3/FS_1/U4_0_2_2  (.A(\mult_20_3/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_20_3/FS_1/P[0][2][2] ),
	.OUT(n3104));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_2  (.A(\mult_20_3/FS_1/PG_int[0][2][2] ),
	.B(\mult_20_3/FS_1/C[1][2][2] ),
	.OUT(N141));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_2  (.A(\mult_20_3/FS_1/G_n_int[0][2][2] ),
	.B(\mult_20_3/FS_1/P[0][2][2] ),
	.OUT(n3103));
   NAND2 \mult_20_3/FS_1/U2_0_2_2  (.A(\mult_20_3/A1[10] ),
	.B(\mult_20_3/A2[10] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_2  (.A(n3101),
	.B(n3102),
	.OUT(\mult_20_3/FS_1/P[0][2][2] ));
   OAI21 \mult_20_3/FS_1/U6_0_2_1  (.OUT(\mult_20_3/FS_1/C[1][2][1] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][0] ),
	.B(n3100),
	.A(n3123));
   OAI21 \mult_20_3/FS_1/U5_0_2_1  (.OUT(\mult_20_3/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][1] ),
	.B(n3107),
	.A(\mult_20_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_3/FS_1/U4_0_2_1  (.A(\mult_20_3/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_20_3/FS_1/P[0][2][1] ),
	.OUT(n3099));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_1  (.A(\mult_20_3/FS_1/PG_int[0][2][1] ),
	.B(\mult_20_3/FS_1/C[1][2][1] ),
	.OUT(N140));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_1  (.A(\mult_20_3/FS_1/G_n_int[0][2][1] ),
	.B(\mult_20_3/FS_1/P[0][2][1] ),
	.OUT(n3098));
   NAND2 \mult_20_3/FS_1/U2_0_2_1  (.A(\mult_20_3/A1[9] ),
	.B(\mult_20_3/A2[9] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_1  (.A(n3096),
	.B(n3097),
	.OUT(\mult_20_3/FS_1/P[0][2][1] ));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_0  (.A(\mult_20_3/FS_1/PG_int[0][2][0] ),
	.B(\mult_20_3/FS_1/C[1][2][0] ),
	.OUT(N139));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_0  (.A(\mult_20_3/FS_1/G_n_int[0][2][0] ),
	.B(\mult_20_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3095));
   NAND2 \mult_20_3/FS_1/U2_0_2_0  (.A(\mult_20_3/A1[8] ),
	.B(\mult_20_3/A2[8] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_0  (.A(n3093),
	.B(n3094),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_20_3/FS_1/U3_B_0_1_3  (.A(\mult_20_3/FS_1/G_n_int[0][1][3] ),
	.B(\mult_20_3/FS_1/P[0][1][3] ),
	.OUT(n3092));
   NAND2 \mult_20_3/FS_1/U2_0_1_3  (.A(\mult_20_3/A1[7] ),
	.B(\mult_20_3/A2[7] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_20_3/FS_1/U1_0_1_3  (.A(n3090),
	.B(n3091),
	.OUT(\mult_20_3/FS_1/P[0][1][3] ));
   inverter \mult_20_3/AN1_7  (.IN(matrix12[7]),
	.OUT(\mult_20_3/A_not[7] ));
   inverter \mult_20_3/AN1_6  (.IN(matrix12[6]),
	.OUT(\mult_20_3/A_notx [6]));
   inverter \mult_20_3/AN1_5  (.IN(matrix12[5]),
	.OUT(\mult_20_3/A_notx [5]));
   inverter \mult_20_3/AN1_4  (.IN(matrix12[4]),
	.OUT(\mult_20_3/A_notx [4]));
   inverter \mult_20_3/AN1_3  (.IN(matrix12[3]),
	.OUT(\mult_20_3/A_notx [3]));
   inverter \mult_20_3/AN1_2  (.IN(matrix12[2]),
	.OUT(\mult_20_3/A_notx [2]));
   inverter \mult_20_3/AN1_1  (.IN(matrix12[1]),
	.OUT(\mult_20_3/A_notx [1]));
   inverter \mult_20_3/AN1_0  (.IN(matrix12[0]),
	.OUT(\mult_20_3/A_notx [0]));
   inverter \mult_20_3/AN1_7_0  (.IN(vector_2[7]),
	.OUT(\mult_20_3/B_not[7] ));
   inverter \mult_20_3/AN1_6_0  (.IN(vector_2[6]),
	.OUT(\mult_20_3/B_notx [6]));
   inverter \mult_20_3/AN1_5_0  (.IN(vector_2[5]),
	.OUT(\mult_20_3/B_notx [5]));
   inverter \mult_20_3/AN1_4_0  (.IN(vector_2[4]),
	.OUT(\mult_20_3/B_notx [4]));
   inverter \mult_20_3/AN1_3_0  (.IN(vector_2[3]),
	.OUT(\mult_20_3/B_notx [3]));
   inverter \mult_20_3/AN1_2_0  (.IN(vector_2[2]),
	.OUT(\mult_20_3/B_notx [2]));
   inverter \mult_20_3/AN1_1_0  (.IN(vector_2[1]),
	.OUT(\mult_20_3/B_notx [1]));
   inverter \mult_20_3/AN1_0_0  (.IN(vector_2[0]),
	.OUT(\mult_20_3/B_notx [0]));
   NOR2 \mult_20_3/AN1_7_7  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[7][7] ));
   NOR2 \mult_20_3/AN3_7_6  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[7][6] ));
   NOR2 \mult_20_3/AN3_7_5  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[7][5] ));
   NOR2 \mult_20_3/AN3_7_4  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[7][4] ));
   NOR2 \mult_20_3/AN3_7_3  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[7][3] ));
   NOR2 \mult_20_3/AN3_7_2  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[7][2] ));
   NOR2 \mult_20_3/AN3_7_1  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[7][1] ));
   NOR2 \mult_20_3/AN3_7_0  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[7][0] ));
   NOR2 \mult_20_3/AN2_6_7  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[6][7] ));
   NOR2 \mult_20_3/AN1_6_6  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[6][6] ));
   NOR2 \mult_20_3/AN1_6_5  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[6][5] ));
   NOR2 \mult_20_3/AN1_6_4  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[6][4] ));
   NOR2 \mult_20_3/AN1_6_3  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[6][3] ));
   NOR2 \mult_20_3/AN1_6_2  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[6][2] ));
   NOR2 \mult_20_3/AN1_6_1  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[6][1] ));
   NOR2 \mult_20_3/AN1_6_0_0  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[6][0] ));
   NOR2 \mult_20_3/AN2_5_7  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[5][7] ));
   NOR2 \mult_20_3/AN1_5_6  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[5][6] ));
   NOR2 \mult_20_3/AN1_5_5  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[5][5] ));
   NOR2 \mult_20_3/AN1_5_4  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[5][4] ));
   NOR2 \mult_20_3/AN1_5_3  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[5][3] ));
   NOR2 \mult_20_3/AN1_5_2  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[5][2] ));
   NOR2 \mult_20_3/AN1_5_1  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[5][1] ));
   NOR2 \mult_20_3/AN1_5_0_0  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[5][0] ));
   NOR2 \mult_20_3/AN2_4_7  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[4][7] ));
   NOR2 \mult_20_3/AN1_4_6  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[4][6] ));
   NOR2 \mult_20_3/AN1_4_5  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[4][5] ));
   NOR2 \mult_20_3/AN1_4_4  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[4][4] ));
   NOR2 \mult_20_3/AN1_4_3  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[4][3] ));
   NOR2 \mult_20_3/AN1_4_2  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[4][2] ));
   NOR2 \mult_20_3/AN1_4_1  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[4][1] ));
   NOR2 \mult_20_3/AN1_4_0_0  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[4][0] ));
   NOR2 \mult_20_3/AN2_3_7  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[3][7] ));
   NOR2 \mult_20_3/AN1_3_6  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[3][6] ));
   NOR2 \mult_20_3/AN1_3_5  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[3][5] ));
   NOR2 \mult_20_3/AN1_3_4  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[3][4] ));
   NOR2 \mult_20_3/AN1_3_3  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[3][3] ));
   NOR2 \mult_20_3/AN1_3_2  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[3][2] ));
   NOR2 \mult_20_3/AN1_3_1  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[3][1] ));
   NOR2 \mult_20_3/AN1_3_0_0  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[3][0] ));
   NOR2 \mult_20_3/AN2_2_7  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[2][7] ));
   NOR2 \mult_20_3/AN1_2_6  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[2][6] ));
   NOR2 \mult_20_3/AN1_2_5  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[2][5] ));
   NOR2 \mult_20_3/AN1_2_4  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[2][4] ));
   NOR2 \mult_20_3/AN1_2_3  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[2][3] ));
   NOR2 \mult_20_3/AN1_2_2  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[2][2] ));
   NOR2 \mult_20_3/AN1_2_1  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[2][1] ));
   NOR2 \mult_20_3/AN1_2_0_0  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[2][0] ));
   NOR2 \mult_20_3/AN2_1_7  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[1][7] ));
   NOR2 \mult_20_3/AN1_1_6  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[1][6] ));
   NOR2 \mult_20_3/AN1_1_5  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[1][5] ));
   NOR2 \mult_20_3/AN1_1_4  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[1][4] ));
   NOR2 \mult_20_3/AN1_1_3  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[1][3] ));
   NOR2 \mult_20_3/AN1_1_2  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[1][2] ));
   NOR2 \mult_20_3/AN1_1_1  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[1][1] ));
   NOR2 \mult_20_3/AN1_1_0_0  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[1][0] ));
   NOR2 \mult_20_3/AN2_0_7  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[0][7] ));
   NOR2 \mult_20_3/AN1_0_6  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[0][6] ));
   NOR2 \mult_20_3/AN1_0_5  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[0][5] ));
   NOR2 \mult_20_3/AN1_0_4  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[0][4] ));
   NOR2 \mult_20_3/AN1_0_3  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[0][3] ));
   NOR2 \mult_20_3/AN1_0_2  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[0][2] ));
   NOR2 \mult_20_3/AN1_0_1  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[0][1] ));
   NOR2 \mult_20_3/AN1_0_0_0  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(N129));
   OAI21 \mult_20_2/FS_1/U6_1_0_3  (.OUT(\mult_20_2/FS_1/C[1][3][0] ),
	.C(n3075),
	.B(n3074),
	.A(n3073));
   OAI21 \mult_20_2/FS_1/U6_0_3_1  (.OUT(\mult_20_2/FS_1/C[1][3][1] ),
	.C(\mult_20_2/FS_1/G_n_int[0][3][0] ),
	.B(n3071),
	.A(n3070));
   XOR2 \mult_20_2/FS_1/U3_C_0_3_1  (.A(\mult_20_2/FS_1/PG_int[0][3][1] ),
	.B(\mult_20_2/FS_1/C[1][3][1] ),
	.OUT(N112));
   XOR2 \mult_20_2/FS_1/U3_C_0_3_0  (.A(\mult_20_2/FS_1/PG_int[0][3][0] ),
	.B(\mult_20_2/FS_1/C[1][3][0] ),
	.OUT(N111));
   NAND2 \mult_20_2/FS_1/U3_B_0_3_0  (.A(\mult_20_2/FS_1/G_n_int[0][3][0] ),
	.B(\mult_20_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3067));
   NAND2 \mult_20_2/FS_1/U2_0_3_0  (.A(\mult_20_2/A1[12] ),
	.B(\mult_20_2/A2[12] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_20_2/FS_1/U1_0_3_0  (.A(n3065),
	.B(n3066),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_20_2/FS_1/U6_0_2_3  (.OUT(\mult_20_2/FS_1/C[1][2][3] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][2] ),
	.B(n3064),
	.A(n3063));
   OAI21 \mult_20_2/FS_1/U5_0_2_3  (.OUT(\mult_20_2/FS_1/G[1][0][2] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][3] ),
	.B(n3062),
	.A(n3061));
   NAND2 \mult_20_2/FS_1/U4_0_2_3  (.A(\mult_20_2/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_20_2/FS_1/P[0][2][3] ),
	.OUT(n3074));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_3  (.A(\mult_20_2/FS_1/PG_int[0][2][3] ),
	.B(\mult_20_2/FS_1/C[1][2][3] ),
	.OUT(N110));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_3  (.A(\mult_20_2/FS_1/G_n_int[0][2][3] ),
	.B(\mult_20_2/FS_1/P[0][2][3] ),
	.OUT(n3060));
   NAND2 \mult_20_2/FS_1/U2_0_2_3  (.A(\mult_20_2/A1[11] ),
	.B(\mult_20_2/A2[11] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_3  (.A(n3058),
	.B(n3059),
	.OUT(\mult_20_2/FS_1/P[0][2][3] ));
   OAI21 \mult_20_2/FS_1/U6_0_2_2  (.OUT(\mult_20_2/FS_1/C[1][2][2] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][1] ),
	.B(n3057),
	.A(n3056));
   OAI21 \mult_20_2/FS_1/U5_0_2_2  (.OUT(\mult_20_2/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][2] ),
	.B(n3064),
	.A(n3055));
   NAND2 \mult_20_2/FS_1/U4_0_2_2  (.A(\mult_20_2/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_20_2/FS_1/P[0][2][2] ),
	.OUT(n3054));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_2  (.A(\mult_20_2/FS_1/PG_int[0][2][2] ),
	.B(\mult_20_2/FS_1/C[1][2][2] ),
	.OUT(N109));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_2  (.A(\mult_20_2/FS_1/G_n_int[0][2][2] ),
	.B(\mult_20_2/FS_1/P[0][2][2] ),
	.OUT(n3053));
   NAND2 \mult_20_2/FS_1/U2_0_2_2  (.A(\mult_20_2/A1[10] ),
	.B(\mult_20_2/A2[10] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_2  (.A(n3051),
	.B(n3052),
	.OUT(\mult_20_2/FS_1/P[0][2][2] ));
   OAI21 \mult_20_2/FS_1/U6_0_2_1  (.OUT(\mult_20_2/FS_1/C[1][2][1] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][0] ),
	.B(n3050),
	.A(n3073));
   OAI21 \mult_20_2/FS_1/U5_0_2_1  (.OUT(\mult_20_2/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][1] ),
	.B(n3057),
	.A(\mult_20_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_2/FS_1/U4_0_2_1  (.A(\mult_20_2/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_20_2/FS_1/P[0][2][1] ),
	.OUT(n3049));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_1  (.A(\mult_20_2/FS_1/PG_int[0][2][1] ),
	.B(\mult_20_2/FS_1/C[1][2][1] ),
	.OUT(N108));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_1  (.A(\mult_20_2/FS_1/G_n_int[0][2][1] ),
	.B(\mult_20_2/FS_1/P[0][2][1] ),
	.OUT(n3048));
   NAND2 \mult_20_2/FS_1/U2_0_2_1  (.A(\mult_20_2/A1[9] ),
	.B(\mult_20_2/A2[9] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_1  (.A(n3046),
	.B(n3047),
	.OUT(\mult_20_2/FS_1/P[0][2][1] ));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_0  (.A(\mult_20_2/FS_1/PG_int[0][2][0] ),
	.B(\mult_20_2/FS_1/C[1][2][0] ),
	.OUT(N107));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_0  (.A(\mult_20_2/FS_1/G_n_int[0][2][0] ),
	.B(\mult_20_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3045));
   NAND2 \mult_20_2/FS_1/U2_0_2_0  (.A(\mult_20_2/A1[8] ),
	.B(\mult_20_2/A2[8] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_0  (.A(n3043),
	.B(n3044),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_20_2/FS_1/U3_B_0_1_3  (.A(\mult_20_2/FS_1/G_n_int[0][1][3] ),
	.B(\mult_20_2/FS_1/P[0][1][3] ),
	.OUT(n3042));
   NAND2 \mult_20_2/FS_1/U2_0_1_3  (.A(\mult_20_2/A1[7] ),
	.B(\mult_20_2/A2[7] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_20_2/FS_1/U1_0_1_3  (.A(n3040),
	.B(n3041),
	.OUT(\mult_20_2/FS_1/P[0][1][3] ));
   inverter \mult_20_2/AN1_7  (.IN(matrix11[7]),
	.OUT(\mult_20_2/A_not[7] ));
   inverter \mult_20_2/AN1_6  (.IN(matrix11[6]),
	.OUT(\mult_20_2/A_notx [6]));
   inverter \mult_20_2/AN1_5  (.IN(matrix11[5]),
	.OUT(\mult_20_2/A_notx [5]));
   inverter \mult_20_2/AN1_4  (.IN(matrix11[4]),
	.OUT(\mult_20_2/A_notx [4]));
   inverter \mult_20_2/AN1_3  (.IN(matrix11[3]),
	.OUT(\mult_20_2/A_notx [3]));
   inverter \mult_20_2/AN1_2  (.IN(matrix11[2]),
	.OUT(\mult_20_2/A_notx [2]));
   inverter \mult_20_2/AN1_1  (.IN(matrix11[1]),
	.OUT(\mult_20_2/A_notx [1]));
   inverter \mult_20_2/AN1_0  (.IN(matrix11[0]),
	.OUT(\mult_20_2/A_notx [0]));
   inverter \mult_20_2/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_20_2/B_not[7] ));
   inverter \mult_20_2/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_20_2/B_notx [6]));
   inverter \mult_20_2/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_20_2/B_notx [5]));
   inverter \mult_20_2/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_20_2/B_notx [4]));
   inverter \mult_20_2/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_20_2/B_notx [3]));
   inverter \mult_20_2/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_20_2/B_notx [2]));
   inverter \mult_20_2/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_20_2/B_notx [1]));
   inverter \mult_20_2/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_20_2/B_notx [0]));
   NOR2 \mult_20_2/AN1_7_7  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[7][7] ));
   NOR2 \mult_20_2/AN3_7_6  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[7][6] ));
   NOR2 \mult_20_2/AN3_7_5  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[7][5] ));
   NOR2 \mult_20_2/AN3_7_4  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[7][4] ));
   NOR2 \mult_20_2/AN3_7_3  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[7][3] ));
   NOR2 \mult_20_2/AN3_7_2  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[7][2] ));
   NOR2 \mult_20_2/AN3_7_1  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[7][1] ));
   NOR2 \mult_20_2/AN3_7_0  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[7][0] ));
   NOR2 \mult_20_2/AN2_6_7  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[6][7] ));
   NOR2 \mult_20_2/AN1_6_6  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[6][6] ));
   NOR2 \mult_20_2/AN1_6_5  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[6][5] ));
   NOR2 \mult_20_2/AN1_6_4  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[6][4] ));
   NOR2 \mult_20_2/AN1_6_3  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[6][3] ));
   NOR2 \mult_20_2/AN1_6_2  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[6][2] ));
   NOR2 \mult_20_2/AN1_6_1  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[6][1] ));
   NOR2 \mult_20_2/AN1_6_0_0  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[6][0] ));
   NOR2 \mult_20_2/AN2_5_7  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[5][7] ));
   NOR2 \mult_20_2/AN1_5_6  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[5][6] ));
   NOR2 \mult_20_2/AN1_5_5  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[5][5] ));
   NOR2 \mult_20_2/AN1_5_4  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[5][4] ));
   NOR2 \mult_20_2/AN1_5_3  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[5][3] ));
   NOR2 \mult_20_2/AN1_5_2  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[5][2] ));
   NOR2 \mult_20_2/AN1_5_1  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[5][1] ));
   NOR2 \mult_20_2/AN1_5_0_0  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[5][0] ));
   NOR2 \mult_20_2/AN2_4_7  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[4][7] ));
   NOR2 \mult_20_2/AN1_4_6  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[4][6] ));
   NOR2 \mult_20_2/AN1_4_5  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[4][5] ));
   NOR2 \mult_20_2/AN1_4_4  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[4][4] ));
   NOR2 \mult_20_2/AN1_4_3  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[4][3] ));
   NOR2 \mult_20_2/AN1_4_2  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[4][2] ));
   NOR2 \mult_20_2/AN1_4_1  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[4][1] ));
   NOR2 \mult_20_2/AN1_4_0_0  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[4][0] ));
   NOR2 \mult_20_2/AN2_3_7  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[3][7] ));
   NOR2 \mult_20_2/AN1_3_6  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[3][6] ));
   NOR2 \mult_20_2/AN1_3_5  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[3][5] ));
   NOR2 \mult_20_2/AN1_3_4  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[3][4] ));
   NOR2 \mult_20_2/AN1_3_3  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[3][3] ));
   NOR2 \mult_20_2/AN1_3_2  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[3][2] ));
   NOR2 \mult_20_2/AN1_3_1  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[3][1] ));
   NOR2 \mult_20_2/AN1_3_0_0  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[3][0] ));
   NOR2 \mult_20_2/AN2_2_7  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[2][7] ));
   NOR2 \mult_20_2/AN1_2_6  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[2][6] ));
   NOR2 \mult_20_2/AN1_2_5  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[2][5] ));
   NOR2 \mult_20_2/AN1_2_4  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[2][4] ));
   NOR2 \mult_20_2/AN1_2_3  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[2][3] ));
   NOR2 \mult_20_2/AN1_2_2  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[2][2] ));
   NOR2 \mult_20_2/AN1_2_1  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[2][1] ));
   NOR2 \mult_20_2/AN1_2_0_0  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[2][0] ));
   NOR2 \mult_20_2/AN2_1_7  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[1][7] ));
   NOR2 \mult_20_2/AN1_1_6  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[1][6] ));
   NOR2 \mult_20_2/AN1_1_5  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[1][5] ));
   NOR2 \mult_20_2/AN1_1_4  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[1][4] ));
   NOR2 \mult_20_2/AN1_1_3  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[1][3] ));
   NOR2 \mult_20_2/AN1_1_2  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[1][2] ));
   NOR2 \mult_20_2/AN1_1_1  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[1][1] ));
   NOR2 \mult_20_2/AN1_1_0_0  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[1][0] ));
   NOR2 \mult_20_2/AN2_0_7  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[0][7] ));
   NOR2 \mult_20_2/AN1_0_6  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[0][6] ));
   NOR2 \mult_20_2/AN1_0_5  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[0][5] ));
   NOR2 \mult_20_2/AN1_0_4  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[0][4] ));
   NOR2 \mult_20_2/AN1_0_3  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[0][3] ));
   NOR2 \mult_20_2/AN1_0_2  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[0][2] ));
   NOR2 \mult_20_2/AN1_0_1  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[0][1] ));
   NOR2 \mult_20_2/AN1_0_0_0  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(N97));
   OAI21 \mult_20/FS_1/U6_1_0_3  (.OUT(\mult_20/FS_1/C[1][3][0] ),
	.C(n3025),
	.B(n3024),
	.A(n3023));
   OAI21 \mult_20/FS_1/U6_0_3_1  (.OUT(\mult_20/FS_1/C[1][3][1] ),
	.C(\mult_20/FS_1/G_n_int[0][3][0] ),
	.B(n3021),
	.A(n3020));
   XOR2 \mult_20/FS_1/U3_C_0_3_1  (.A(\mult_20/FS_1/PG_int[0][3][1] ),
	.B(\mult_20/FS_1/C[1][3][1] ),
	.OUT(N96));
   XOR2 \mult_20/FS_1/U3_C_0_3_0  (.A(\mult_20/FS_1/PG_int[0][3][0] ),
	.B(\mult_20/FS_1/C[1][3][0] ),
	.OUT(N95));
   NAND2 \mult_20/FS_1/U3_B_0_3_0  (.A(\mult_20/FS_1/G_n_int[0][3][0] ),
	.B(\mult_20/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3017));
   NAND2 \mult_20/FS_1/U2_0_3_0  (.A(\mult_20/A1[12] ),
	.B(\mult_20/A2[12] ),
	.OUT(\mult_20/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_20/FS_1/U1_0_3_0  (.A(n3015),
	.B(n3016),
	.OUT(\mult_20/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_20/FS_1/U6_0_2_3  (.OUT(\mult_20/FS_1/C[1][2][3] ),
	.C(\mult_20/FS_1/G_n_int[0][2][2] ),
	.B(n3014),
	.A(n3013));
   OAI21 \mult_20/FS_1/U5_0_2_3  (.OUT(\mult_20/FS_1/G[1][0][2] ),
	.C(\mult_20/FS_1/G_n_int[0][2][3] ),
	.B(n3012),
	.A(n3011));
   NAND2 \mult_20/FS_1/U4_0_2_3  (.A(\mult_20/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_20/FS_1/P[0][2][3] ),
	.OUT(n3024));
   XOR2 \mult_20/FS_1/U3_C_0_2_3  (.A(\mult_20/FS_1/PG_int[0][2][3] ),
	.B(\mult_20/FS_1/C[1][2][3] ),
	.OUT(N94));
   NAND2 \mult_20/FS_1/U3_B_0_2_3  (.A(\mult_20/FS_1/G_n_int[0][2][3] ),
	.B(\mult_20/FS_1/P[0][2][3] ),
	.OUT(n3010));
   NAND2 \mult_20/FS_1/U2_0_2_3  (.A(\mult_20/A1[11] ),
	.B(\mult_20/A2[11] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_20/FS_1/U1_0_2_3  (.A(n3008),
	.B(n3009),
	.OUT(\mult_20/FS_1/P[0][2][3] ));
   OAI21 \mult_20/FS_1/U6_0_2_2  (.OUT(\mult_20/FS_1/C[1][2][2] ),
	.C(\mult_20/FS_1/G_n_int[0][2][1] ),
	.B(n3007),
	.A(n3006));
   OAI21 \mult_20/FS_1/U5_0_2_2  (.OUT(\mult_20/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_20/FS_1/G_n_int[0][2][2] ),
	.B(n3014),
	.A(n3005));
   NAND2 \mult_20/FS_1/U4_0_2_2  (.A(\mult_20/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_20/FS_1/P[0][2][2] ),
	.OUT(n3004));
   XOR2 \mult_20/FS_1/U3_C_0_2_2  (.A(\mult_20/FS_1/PG_int[0][2][2] ),
	.B(\mult_20/FS_1/C[1][2][2] ),
	.OUT(N93));
   NAND2 \mult_20/FS_1/U3_B_0_2_2  (.A(\mult_20/FS_1/G_n_int[0][2][2] ),
	.B(\mult_20/FS_1/P[0][2][2] ),
	.OUT(n3003));
   NAND2 \mult_20/FS_1/U2_0_2_2  (.A(\mult_20/A1[10] ),
	.B(\mult_20/A2[10] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_20/FS_1/U1_0_2_2  (.A(n3001),
	.B(n3002),
	.OUT(\mult_20/FS_1/P[0][2][2] ));
   OAI21 \mult_20/FS_1/U6_0_2_1  (.OUT(\mult_20/FS_1/C[1][2][1] ),
	.C(\mult_20/FS_1/G_n_int[0][2][0] ),
	.B(n3000),
	.A(n3023));
   OAI21 \mult_20/FS_1/U5_0_2_1  (.OUT(\mult_20/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_20/FS_1/G_n_int[0][2][1] ),
	.B(n3007),
	.A(\mult_20/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20/FS_1/U4_0_2_1  (.A(\mult_20/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_20/FS_1/P[0][2][1] ),
	.OUT(n2999));
   XOR2 \mult_20/FS_1/U3_C_0_2_1  (.A(\mult_20/FS_1/PG_int[0][2][1] ),
	.B(\mult_20/FS_1/C[1][2][1] ),
	.OUT(N92));
   NAND2 \mult_20/FS_1/U3_B_0_2_1  (.A(\mult_20/FS_1/G_n_int[0][2][1] ),
	.B(\mult_20/FS_1/P[0][2][1] ),
	.OUT(n2998));
   NAND2 \mult_20/FS_1/U2_0_2_1  (.A(\mult_20/A1[9] ),
	.B(\mult_20/A2[9] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_20/FS_1/U1_0_2_1  (.A(n2996),
	.B(n2997),
	.OUT(\mult_20/FS_1/P[0][2][1] ));
   XOR2 \mult_20/FS_1/U3_C_0_2_0  (.A(\mult_20/FS_1/PG_int[0][2][0] ),
	.B(\mult_20/FS_1/C[1][2][0] ),
	.OUT(N91));
   NAND2 \mult_20/FS_1/U3_B_0_2_0  (.A(\mult_20/FS_1/G_n_int[0][2][0] ),
	.B(\mult_20/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2995));
   NAND2 \mult_20/FS_1/U2_0_2_0  (.A(\mult_20/A1[8] ),
	.B(\mult_20/A2[8] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20/FS_1/U1_0_2_0  (.A(n2993),
	.B(n2994),
	.OUT(\mult_20/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_20/FS_1/U3_B_0_1_3  (.A(\mult_20/FS_1/G_n_int[0][1][3] ),
	.B(\mult_20/FS_1/P[0][1][3] ),
	.OUT(n2992));
   NAND2 \mult_20/FS_1/U2_0_1_3  (.A(\mult_20/A1[7] ),
	.B(\mult_20/A2[7] ),
	.OUT(\mult_20/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_20/FS_1/U1_0_1_3  (.A(n2990),
	.B(n2991),
	.OUT(\mult_20/FS_1/P[0][1][3] ));
   inverter \mult_20/AN1_7  (.IN(matrix10[7]),
	.OUT(\mult_20/A_not[7] ));
   inverter \mult_20/AN1_6  (.IN(matrix10[6]),
	.OUT(\mult_20/A_notx [6]));
   inverter \mult_20/AN1_5  (.IN(matrix10[5]),
	.OUT(\mult_20/A_notx [5]));
   inverter \mult_20/AN1_4  (.IN(matrix10[4]),
	.OUT(\mult_20/A_notx [4]));
   inverter \mult_20/AN1_3  (.IN(matrix10[3]),
	.OUT(\mult_20/A_notx [3]));
   inverter \mult_20/AN1_2  (.IN(matrix10[2]),
	.OUT(\mult_20/A_notx [2]));
   inverter \mult_20/AN1_1  (.IN(matrix10[1]),
	.OUT(\mult_20/A_notx [1]));
   inverter \mult_20/AN1_0  (.IN(matrix10[0]),
	.OUT(\mult_20/A_notx [0]));
   inverter \mult_20/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_20/B_not[7] ));
   inverter \mult_20/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_20/B_notx [6]));
   inverter \mult_20/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_20/B_notx [5]));
   inverter \mult_20/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_20/B_notx [4]));
   inverter \mult_20/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_20/B_notx [3]));
   inverter \mult_20/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_20/B_notx [2]));
   inverter \mult_20/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_20/B_notx [1]));
   inverter \mult_20/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_20/B_notx [0]));
   NOR2 \mult_20/AN1_7_7  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[7][7] ));
   NOR2 \mult_20/AN3_7_6  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[7][6] ));
   NOR2 \mult_20/AN3_7_5  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[7][5] ));
   NOR2 \mult_20/AN3_7_4  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[7][4] ));
   NOR2 \mult_20/AN3_7_3  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[7][3] ));
   NOR2 \mult_20/AN3_7_2  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[7][2] ));
   NOR2 \mult_20/AN3_7_1  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[7][1] ));
   NOR2 \mult_20/AN3_7_0  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[7][0] ));
   NOR2 \mult_20/AN2_6_7  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[6][7] ));
   NOR2 \mult_20/AN1_6_6  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[6][6] ));
   NOR2 \mult_20/AN1_6_5  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[6][5] ));
   NOR2 \mult_20/AN1_6_4  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[6][4] ));
   NOR2 \mult_20/AN1_6_3  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[6][3] ));
   NOR2 \mult_20/AN1_6_2  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[6][2] ));
   NOR2 \mult_20/AN1_6_1  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[6][1] ));
   NOR2 \mult_20/AN1_6_0_0  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[6][0] ));
   NOR2 \mult_20/AN2_5_7  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[5][7] ));
   NOR2 \mult_20/AN1_5_6  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[5][6] ));
   NOR2 \mult_20/AN1_5_5  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[5][5] ));
   NOR2 \mult_20/AN1_5_4  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[5][4] ));
   NOR2 \mult_20/AN1_5_3  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[5][3] ));
   NOR2 \mult_20/AN1_5_2  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[5][2] ));
   NOR2 \mult_20/AN1_5_1  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[5][1] ));
   NOR2 \mult_20/AN1_5_0_0  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[5][0] ));
   NOR2 \mult_20/AN2_4_7  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[4][7] ));
   NOR2 \mult_20/AN1_4_6  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[4][6] ));
   NOR2 \mult_20/AN1_4_5  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[4][5] ));
   NOR2 \mult_20/AN1_4_4  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[4][4] ));
   NOR2 \mult_20/AN1_4_3  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[4][3] ));
   NOR2 \mult_20/AN1_4_2  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[4][2] ));
   NOR2 \mult_20/AN1_4_1  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[4][1] ));
   NOR2 \mult_20/AN1_4_0_0  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[4][0] ));
   NOR2 \mult_20/AN2_3_7  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[3][7] ));
   NOR2 \mult_20/AN1_3_6  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[3][6] ));
   NOR2 \mult_20/AN1_3_5  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[3][5] ));
   NOR2 \mult_20/AN1_3_4  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[3][4] ));
   NOR2 \mult_20/AN1_3_3  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[3][3] ));
   NOR2 \mult_20/AN1_3_2  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[3][2] ));
   NOR2 \mult_20/AN1_3_1  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[3][1] ));
   NOR2 \mult_20/AN1_3_0_0  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[3][0] ));
   NOR2 \mult_20/AN2_2_7  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[2][7] ));
   NOR2 \mult_20/AN1_2_6  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[2][6] ));
   NOR2 \mult_20/AN1_2_5  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[2][5] ));
   NOR2 \mult_20/AN1_2_4  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[2][4] ));
   NOR2 \mult_20/AN1_2_3  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[2][3] ));
   NOR2 \mult_20/AN1_2_2  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[2][2] ));
   NOR2 \mult_20/AN1_2_1  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[2][1] ));
   NOR2 \mult_20/AN1_2_0_0  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[2][0] ));
   NOR2 \mult_20/AN2_1_7  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[1][7] ));
   NOR2 \mult_20/AN1_1_6  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[1][6] ));
   NOR2 \mult_20/AN1_1_5  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[1][5] ));
   NOR2 \mult_20/AN1_1_4  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[1][4] ));
   NOR2 \mult_20/AN1_1_3  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[1][3] ));
   NOR2 \mult_20/AN1_1_2  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[1][2] ));
   NOR2 \mult_20/AN1_1_1  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[1][1] ));
   NOR2 \mult_20/AN1_1_0_0  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[1][0] ));
   NOR2 \mult_20/AN2_0_7  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[0][7] ));
   NOR2 \mult_20/AN1_0_6  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[0][6] ));
   NOR2 \mult_20/AN1_0_5  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[0][5] ));
   NOR2 \mult_20/AN1_0_4  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[0][4] ));
   NOR2 \mult_20/AN1_0_3  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[0][3] ));
   NOR2 \mult_20/AN1_0_2  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[0][2] ));
   NOR2 \mult_20/AN1_0_1  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[0][1] ));
   NOR2 \mult_20/AN1_0_0_0  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [0]),
	.OUT(N81));
   OAI21 \mult_19_3/FS_1/U6_1_0_3  (.OUT(\mult_19_3/FS_1/C[1][3][0] ),
	.C(n2975),
	.B(n2974),
	.A(n2973));
   OAI21 \mult_19_3/FS_1/U6_0_3_1  (.OUT(\mult_19_3/FS_1/C[1][3][1] ),
	.C(\mult_19_3/FS_1/G_n_int[0][3][0] ),
	.B(n2971),
	.A(n2970));
   XOR2 \mult_19_3/FS_1/U3_C_0_3_1  (.A(\mult_19_3/FS_1/PG_int[0][3][1] ),
	.B(\mult_19_3/FS_1/C[1][3][1] ),
	.OUT(N64));
   XOR2 \mult_19_3/FS_1/U3_C_0_3_0  (.A(\mult_19_3/FS_1/PG_int[0][3][0] ),
	.B(\mult_19_3/FS_1/C[1][3][0] ),
	.OUT(N63));
   NAND2 \mult_19_3/FS_1/U3_B_0_3_0  (.A(\mult_19_3/FS_1/G_n_int[0][3][0] ),
	.B(\mult_19_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2967));
   NAND2 \mult_19_3/FS_1/U2_0_3_0  (.A(\mult_19_3/A1[12] ),
	.B(\mult_19_3/A2[12] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_19_3/FS_1/U1_0_3_0  (.A(n2965),
	.B(n2966),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_19_3/FS_1/U6_0_2_3  (.OUT(\mult_19_3/FS_1/C[1][2][3] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][2] ),
	.B(n2964),
	.A(n2963));
   OAI21 \mult_19_3/FS_1/U5_0_2_3  (.OUT(\mult_19_3/FS_1/G[1][0][2] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][3] ),
	.B(n2962),
	.A(n2961));
   NAND2 \mult_19_3/FS_1/U4_0_2_3  (.A(\mult_19_3/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_19_3/FS_1/P[0][2][3] ),
	.OUT(n2974));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_3  (.A(\mult_19_3/FS_1/PG_int[0][2][3] ),
	.B(\mult_19_3/FS_1/C[1][2][3] ),
	.OUT(N62));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_3  (.A(\mult_19_3/FS_1/G_n_int[0][2][3] ),
	.B(\mult_19_3/FS_1/P[0][2][3] ),
	.OUT(n2960));
   NAND2 \mult_19_3/FS_1/U2_0_2_3  (.A(\mult_19_3/A1[11] ),
	.B(\mult_19_3/A2[11] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_3  (.A(n2958),
	.B(n2959),
	.OUT(\mult_19_3/FS_1/P[0][2][3] ));
   OAI21 \mult_19_3/FS_1/U6_0_2_2  (.OUT(\mult_19_3/FS_1/C[1][2][2] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][1] ),
	.B(n2957),
	.A(n2956));
   OAI21 \mult_19_3/FS_1/U5_0_2_2  (.OUT(\mult_19_3/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][2] ),
	.B(n2964),
	.A(n2955));
   NAND2 \mult_19_3/FS_1/U4_0_2_2  (.A(\mult_19_3/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_19_3/FS_1/P[0][2][2] ),
	.OUT(n2954));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_2  (.A(\mult_19_3/FS_1/PG_int[0][2][2] ),
	.B(\mult_19_3/FS_1/C[1][2][2] ),
	.OUT(N61));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_2  (.A(\mult_19_3/FS_1/G_n_int[0][2][2] ),
	.B(\mult_19_3/FS_1/P[0][2][2] ),
	.OUT(n2953));
   NAND2 \mult_19_3/FS_1/U2_0_2_2  (.A(\mult_19_3/A1[10] ),
	.B(\mult_19_3/A2[10] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_2  (.A(n2951),
	.B(n2952),
	.OUT(\mult_19_3/FS_1/P[0][2][2] ));
   OAI21 \mult_19_3/FS_1/U6_0_2_1  (.OUT(\mult_19_3/FS_1/C[1][2][1] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][0] ),
	.B(n2950),
	.A(n2973));
   OAI21 \mult_19_3/FS_1/U5_0_2_1  (.OUT(\mult_19_3/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][1] ),
	.B(n2957),
	.A(\mult_19_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_3/FS_1/U4_0_2_1  (.A(\mult_19_3/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_19_3/FS_1/P[0][2][1] ),
	.OUT(n2949));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_1  (.A(\mult_19_3/FS_1/PG_int[0][2][1] ),
	.B(\mult_19_3/FS_1/C[1][2][1] ),
	.OUT(N60));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_1  (.A(\mult_19_3/FS_1/G_n_int[0][2][1] ),
	.B(\mult_19_3/FS_1/P[0][2][1] ),
	.OUT(n2948));
   NAND2 \mult_19_3/FS_1/U2_0_2_1  (.A(\mult_19_3/A1[9] ),
	.B(\mult_19_3/A2[9] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_1  (.A(n2946),
	.B(n2947),
	.OUT(\mult_19_3/FS_1/P[0][2][1] ));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_0  (.A(\mult_19_3/FS_1/PG_int[0][2][0] ),
	.B(\mult_19_3/FS_1/C[1][2][0] ),
	.OUT(N59));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_0  (.A(\mult_19_3/FS_1/G_n_int[0][2][0] ),
	.B(\mult_19_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2945));
   NAND2 \mult_19_3/FS_1/U2_0_2_0  (.A(\mult_19_3/A1[8] ),
	.B(\mult_19_3/A2[8] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_0  (.A(n2943),
	.B(n2944),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_19_3/FS_1/U3_B_0_1_3  (.A(\mult_19_3/FS_1/G_n_int[0][1][3] ),
	.B(\mult_19_3/FS_1/P[0][1][3] ),
	.OUT(n2942));
   NAND2 \mult_19_3/FS_1/U2_0_1_3  (.A(\mult_19_3/A1[7] ),
	.B(\mult_19_3/A2[7] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_19_3/FS_1/U1_0_1_3  (.A(n2940),
	.B(n2941),
	.OUT(\mult_19_3/FS_1/P[0][1][3] ));
   inverter \mult_19_3/AN1_7  (.IN(matrix02[7]),
	.OUT(\mult_19_3/A_not[7] ));
   inverter \mult_19_3/AN1_6  (.IN(matrix02[6]),
	.OUT(\mult_19_3/A_notx [6]));
   inverter \mult_19_3/AN1_5  (.IN(matrix02[5]),
	.OUT(\mult_19_3/A_notx [5]));
   inverter \mult_19_3/AN1_4  (.IN(matrix02[4]),
	.OUT(\mult_19_3/A_notx [4]));
   inverter \mult_19_3/AN1_3  (.IN(matrix02[3]),
	.OUT(\mult_19_3/A_notx [3]));
   inverter \mult_19_3/AN1_2  (.IN(matrix02[2]),
	.OUT(\mult_19_3/A_notx [2]));
   inverter \mult_19_3/AN1_1  (.IN(matrix02[1]),
	.OUT(\mult_19_3/A_notx [1]));
   inverter \mult_19_3/AN1_0  (.IN(matrix02[0]),
	.OUT(\mult_19_3/A_notx [0]));
   inverter \mult_19_3/AN1_7_0  (.IN(vector_2[7]),
	.OUT(\mult_19_3/B_not[7] ));
   inverter \mult_19_3/AN1_6_0  (.IN(vector_2[6]),
	.OUT(\mult_19_3/B_notx [6]));
   inverter \mult_19_3/AN1_5_0  (.IN(vector_2[5]),
	.OUT(\mult_19_3/B_notx [5]));
   inverter \mult_19_3/AN1_4_0  (.IN(vector_2[4]),
	.OUT(\mult_19_3/B_notx [4]));
   inverter \mult_19_3/AN1_3_0  (.IN(vector_2[3]),
	.OUT(\mult_19_3/B_notx [3]));
   inverter \mult_19_3/AN1_2_0  (.IN(vector_2[2]),
	.OUT(\mult_19_3/B_notx [2]));
   inverter \mult_19_3/AN1_1_0  (.IN(vector_2[1]),
	.OUT(\mult_19_3/B_notx [1]));
   inverter \mult_19_3/AN1_0_0  (.IN(vector_2[0]),
	.OUT(\mult_19_3/B_notx [0]));
   NOR2 \mult_19_3/AN1_7_7  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[7][7] ));
   NOR2 \mult_19_3/AN3_7_6  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[7][6] ));
   NOR2 \mult_19_3/AN3_7_5  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[7][5] ));
   NOR2 \mult_19_3/AN3_7_4  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[7][4] ));
   NOR2 \mult_19_3/AN3_7_3  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[7][3] ));
   NOR2 \mult_19_3/AN3_7_2  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[7][2] ));
   NOR2 \mult_19_3/AN3_7_1  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[7][1] ));
   NOR2 \mult_19_3/AN3_7_0  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[7][0] ));
   NOR2 \mult_19_3/AN2_6_7  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[6][7] ));
   NOR2 \mult_19_3/AN1_6_6  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[6][6] ));
   NOR2 \mult_19_3/AN1_6_5  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[6][5] ));
   NOR2 \mult_19_3/AN1_6_4  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[6][4] ));
   NOR2 \mult_19_3/AN1_6_3  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[6][3] ));
   NOR2 \mult_19_3/AN1_6_2  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[6][2] ));
   NOR2 \mult_19_3/AN1_6_1  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[6][1] ));
   NOR2 \mult_19_3/AN1_6_0_0  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[6][0] ));
   NOR2 \mult_19_3/AN2_5_7  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[5][7] ));
   NOR2 \mult_19_3/AN1_5_6  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[5][6] ));
   NOR2 \mult_19_3/AN1_5_5  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[5][5] ));
   NOR2 \mult_19_3/AN1_5_4  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[5][4] ));
   NOR2 \mult_19_3/AN1_5_3  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[5][3] ));
   NOR2 \mult_19_3/AN1_5_2  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[5][2] ));
   NOR2 \mult_19_3/AN1_5_1  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[5][1] ));
   NOR2 \mult_19_3/AN1_5_0_0  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[5][0] ));
   NOR2 \mult_19_3/AN2_4_7  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[4][7] ));
   NOR2 \mult_19_3/AN1_4_6  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[4][6] ));
   NOR2 \mult_19_3/AN1_4_5  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[4][5] ));
   NOR2 \mult_19_3/AN1_4_4  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[4][4] ));
   NOR2 \mult_19_3/AN1_4_3  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[4][3] ));
   NOR2 \mult_19_3/AN1_4_2  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[4][2] ));
   NOR2 \mult_19_3/AN1_4_1  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[4][1] ));
   NOR2 \mult_19_3/AN1_4_0_0  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[4][0] ));
   NOR2 \mult_19_3/AN2_3_7  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[3][7] ));
   NOR2 \mult_19_3/AN1_3_6  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[3][6] ));
   NOR2 \mult_19_3/AN1_3_5  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[3][5] ));
   NOR2 \mult_19_3/AN1_3_4  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[3][4] ));
   NOR2 \mult_19_3/AN1_3_3  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[3][3] ));
   NOR2 \mult_19_3/AN1_3_2  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[3][2] ));
   NOR2 \mult_19_3/AN1_3_1  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[3][1] ));
   NOR2 \mult_19_3/AN1_3_0_0  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[3][0] ));
   NOR2 \mult_19_3/AN2_2_7  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[2][7] ));
   NOR2 \mult_19_3/AN1_2_6  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[2][6] ));
   NOR2 \mult_19_3/AN1_2_5  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[2][5] ));
   NOR2 \mult_19_3/AN1_2_4  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[2][4] ));
   NOR2 \mult_19_3/AN1_2_3  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[2][3] ));
   NOR2 \mult_19_3/AN1_2_2  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[2][2] ));
   NOR2 \mult_19_3/AN1_2_1  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[2][1] ));
   NOR2 \mult_19_3/AN1_2_0_0  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[2][0] ));
   NOR2 \mult_19_3/AN2_1_7  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[1][7] ));
   NOR2 \mult_19_3/AN1_1_6  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[1][6] ));
   NOR2 \mult_19_3/AN1_1_5  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[1][5] ));
   NOR2 \mult_19_3/AN1_1_4  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[1][4] ));
   NOR2 \mult_19_3/AN1_1_3  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[1][3] ));
   NOR2 \mult_19_3/AN1_1_2  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[1][2] ));
   NOR2 \mult_19_3/AN1_1_1  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[1][1] ));
   NOR2 \mult_19_3/AN1_1_0_0  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[1][0] ));
   NOR2 \mult_19_3/AN2_0_7  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[0][7] ));
   NOR2 \mult_19_3/AN1_0_6  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[0][6] ));
   NOR2 \mult_19_3/AN1_0_5  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[0][5] ));
   NOR2 \mult_19_3/AN1_0_4  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[0][4] ));
   NOR2 \mult_19_3/AN1_0_3  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[0][3] ));
   NOR2 \mult_19_3/AN1_0_2  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[0][2] ));
   NOR2 \mult_19_3/AN1_0_1  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[0][1] ));
   NOR2 \mult_19_3/AN1_0_0_0  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(N49));
   OAI21 \mult_19_2/FS_1/U6_1_0_3  (.OUT(\mult_19_2/FS_1/C[1][3][0] ),
	.C(n2925),
	.B(n2924),
	.A(n2923));
   OAI21 \mult_19_2/FS_1/U6_0_3_1  (.OUT(\mult_19_2/FS_1/C[1][3][1] ),
	.C(\mult_19_2/FS_1/G_n_int[0][3][0] ),
	.B(n2921),
	.A(n2920));
   XOR2 \mult_19_2/FS_1/U3_C_0_3_1  (.A(\mult_19_2/FS_1/PG_int[0][3][1] ),
	.B(\mult_19_2/FS_1/C[1][3][1] ),
	.OUT(N32));
   XOR2 \mult_19_2/FS_1/U3_C_0_3_0  (.A(\mult_19_2/FS_1/PG_int[0][3][0] ),
	.B(\mult_19_2/FS_1/C[1][3][0] ),
	.OUT(N31));
   NAND2 \mult_19_2/FS_1/U3_B_0_3_0  (.A(\mult_19_2/FS_1/G_n_int[0][3][0] ),
	.B(\mult_19_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2917));
   NAND2 \mult_19_2/FS_1/U2_0_3_0  (.A(\mult_19_2/A1[12] ),
	.B(\mult_19_2/A2[12] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_19_2/FS_1/U1_0_3_0  (.A(n2915),
	.B(n2916),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_19_2/FS_1/U6_0_2_3  (.OUT(\mult_19_2/FS_1/C[1][2][3] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][2] ),
	.B(n2914),
	.A(n2913));
   OAI21 \mult_19_2/FS_1/U5_0_2_3  (.OUT(\mult_19_2/FS_1/G[1][0][2] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][3] ),
	.B(n2912),
	.A(n2911));
   NAND2 \mult_19_2/FS_1/U4_0_2_3  (.A(\mult_19_2/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_19_2/FS_1/P[0][2][3] ),
	.OUT(n2924));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_3  (.A(\mult_19_2/FS_1/PG_int[0][2][3] ),
	.B(\mult_19_2/FS_1/C[1][2][3] ),
	.OUT(N30));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_3  (.A(\mult_19_2/FS_1/G_n_int[0][2][3] ),
	.B(\mult_19_2/FS_1/P[0][2][3] ),
	.OUT(n2910));
   NAND2 \mult_19_2/FS_1/U2_0_2_3  (.A(\mult_19_2/A1[11] ),
	.B(\mult_19_2/A2[11] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_3  (.A(n2908),
	.B(n2909),
	.OUT(\mult_19_2/FS_1/P[0][2][3] ));
   OAI21 \mult_19_2/FS_1/U6_0_2_2  (.OUT(\mult_19_2/FS_1/C[1][2][2] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][1] ),
	.B(n2907),
	.A(n2906));
   OAI21 \mult_19_2/FS_1/U5_0_2_2  (.OUT(\mult_19_2/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][2] ),
	.B(n2914),
	.A(n2905));
   NAND2 \mult_19_2/FS_1/U4_0_2_2  (.A(\mult_19_2/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_19_2/FS_1/P[0][2][2] ),
	.OUT(n2904));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_2  (.A(\mult_19_2/FS_1/PG_int[0][2][2] ),
	.B(\mult_19_2/FS_1/C[1][2][2] ),
	.OUT(N29));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_2  (.A(\mult_19_2/FS_1/G_n_int[0][2][2] ),
	.B(\mult_19_2/FS_1/P[0][2][2] ),
	.OUT(n2903));
   NAND2 \mult_19_2/FS_1/U2_0_2_2  (.A(\mult_19_2/A1[10] ),
	.B(\mult_19_2/A2[10] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_2  (.A(n2901),
	.B(n2902),
	.OUT(\mult_19_2/FS_1/P[0][2][2] ));
   OAI21 \mult_19_2/FS_1/U6_0_2_1  (.OUT(\mult_19_2/FS_1/C[1][2][1] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][0] ),
	.B(n2900),
	.A(n2923));
   OAI21 \mult_19_2/FS_1/U5_0_2_1  (.OUT(\mult_19_2/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][1] ),
	.B(n2907),
	.A(\mult_19_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_2/FS_1/U4_0_2_1  (.A(\mult_19_2/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_19_2/FS_1/P[0][2][1] ),
	.OUT(n2899));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_1  (.A(\mult_19_2/FS_1/PG_int[0][2][1] ),
	.B(\mult_19_2/FS_1/C[1][2][1] ),
	.OUT(N28));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_1  (.A(\mult_19_2/FS_1/G_n_int[0][2][1] ),
	.B(\mult_19_2/FS_1/P[0][2][1] ),
	.OUT(n2898));
   NAND2 \mult_19_2/FS_1/U2_0_2_1  (.A(\mult_19_2/A1[9] ),
	.B(\mult_19_2/A2[9] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_1  (.A(n2896),
	.B(n2897),
	.OUT(\mult_19_2/FS_1/P[0][2][1] ));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_0  (.A(\mult_19_2/FS_1/PG_int[0][2][0] ),
	.B(\mult_19_2/FS_1/C[1][2][0] ),
	.OUT(N27));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_0  (.A(\mult_19_2/FS_1/G_n_int[0][2][0] ),
	.B(\mult_19_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2895));
   NAND2 \mult_19_2/FS_1/U2_0_2_0  (.A(\mult_19_2/A1[8] ),
	.B(\mult_19_2/A2[8] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_0  (.A(n2893),
	.B(n2894),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_19_2/FS_1/U3_B_0_1_3  (.A(\mult_19_2/FS_1/G_n_int[0][1][3] ),
	.B(\mult_19_2/FS_1/P[0][1][3] ),
	.OUT(n2892));
   NAND2 \mult_19_2/FS_1/U2_0_1_3  (.A(\mult_19_2/A1[7] ),
	.B(\mult_19_2/A2[7] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_19_2/FS_1/U1_0_1_3  (.A(n2890),
	.B(n2891),
	.OUT(\mult_19_2/FS_1/P[0][1][3] ));
   inverter \mult_19_2/AN1_7  (.IN(matrix01[7]),
	.OUT(\mult_19_2/A_not[7] ));
   inverter \mult_19_2/AN1_6  (.IN(matrix01[6]),
	.OUT(\mult_19_2/A_notx [6]));
   inverter \mult_19_2/AN1_5  (.IN(matrix01[5]),
	.OUT(\mult_19_2/A_notx [5]));
   inverter \mult_19_2/AN1_4  (.IN(matrix01[4]),
	.OUT(\mult_19_2/A_notx [4]));
   inverter \mult_19_2/AN1_3  (.IN(matrix01[3]),
	.OUT(\mult_19_2/A_notx [3]));
   inverter \mult_19_2/AN1_2  (.IN(matrix01[2]),
	.OUT(\mult_19_2/A_notx [2]));
   inverter \mult_19_2/AN1_1  (.IN(matrix01[1]),
	.OUT(\mult_19_2/A_notx [1]));
   inverter \mult_19_2/AN1_0  (.IN(matrix01[0]),
	.OUT(\mult_19_2/A_notx [0]));
   inverter \mult_19_2/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_19_2/B_not[7] ));
   inverter \mult_19_2/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_19_2/B_notx [6]));
   inverter \mult_19_2/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_19_2/B_notx [5]));
   inverter \mult_19_2/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_19_2/B_notx [4]));
   inverter \mult_19_2/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_19_2/B_notx [3]));
   inverter \mult_19_2/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_19_2/B_notx [2]));
   inverter \mult_19_2/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_19_2/B_notx [1]));
   inverter \mult_19_2/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_19_2/B_notx [0]));
   NOR2 \mult_19_2/AN1_7_7  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[7][7] ));
   NOR2 \mult_19_2/AN3_7_6  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[7][6] ));
   NOR2 \mult_19_2/AN3_7_5  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[7][5] ));
   NOR2 \mult_19_2/AN3_7_4  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[7][4] ));
   NOR2 \mult_19_2/AN3_7_3  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[7][3] ));
   NOR2 \mult_19_2/AN3_7_2  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[7][2] ));
   NOR2 \mult_19_2/AN3_7_1  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[7][1] ));
   NOR2 \mult_19_2/AN3_7_0  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[7][0] ));
   NOR2 \mult_19_2/AN2_6_7  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[6][7] ));
   NOR2 \mult_19_2/AN1_6_6  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[6][6] ));
   NOR2 \mult_19_2/AN1_6_5  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[6][5] ));
   NOR2 \mult_19_2/AN1_6_4  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[6][4] ));
   NOR2 \mult_19_2/AN1_6_3  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[6][3] ));
   NOR2 \mult_19_2/AN1_6_2  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[6][2] ));
   NOR2 \mult_19_2/AN1_6_1  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[6][1] ));
   NOR2 \mult_19_2/AN1_6_0_0  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[6][0] ));
   NOR2 \mult_19_2/AN2_5_7  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[5][7] ));
   NOR2 \mult_19_2/AN1_5_6  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[5][6] ));
   NOR2 \mult_19_2/AN1_5_5  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[5][5] ));
   NOR2 \mult_19_2/AN1_5_4  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[5][4] ));
   NOR2 \mult_19_2/AN1_5_3  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[5][3] ));
   NOR2 \mult_19_2/AN1_5_2  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[5][2] ));
   NOR2 \mult_19_2/AN1_5_1  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[5][1] ));
   NOR2 \mult_19_2/AN1_5_0_0  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[5][0] ));
   NOR2 \mult_19_2/AN2_4_7  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[4][7] ));
   NOR2 \mult_19_2/AN1_4_6  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[4][6] ));
   NOR2 \mult_19_2/AN1_4_5  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[4][5] ));
   NOR2 \mult_19_2/AN1_4_4  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[4][4] ));
   NOR2 \mult_19_2/AN1_4_3  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[4][3] ));
   NOR2 \mult_19_2/AN1_4_2  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[4][2] ));
   NOR2 \mult_19_2/AN1_4_1  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[4][1] ));
   NOR2 \mult_19_2/AN1_4_0_0  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[4][0] ));
   NOR2 \mult_19_2/AN2_3_7  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[3][7] ));
   NOR2 \mult_19_2/AN1_3_6  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[3][6] ));
   NOR2 \mult_19_2/AN1_3_5  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[3][5] ));
   NOR2 \mult_19_2/AN1_3_4  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[3][4] ));
   NOR2 \mult_19_2/AN1_3_3  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[3][3] ));
   NOR2 \mult_19_2/AN1_3_2  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[3][2] ));
   NOR2 \mult_19_2/AN1_3_1  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[3][1] ));
   NOR2 \mult_19_2/AN1_3_0_0  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[3][0] ));
   NOR2 \mult_19_2/AN2_2_7  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[2][7] ));
   NOR2 \mult_19_2/AN1_2_6  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[2][6] ));
   NOR2 \mult_19_2/AN1_2_5  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[2][5] ));
   NOR2 \mult_19_2/AN1_2_4  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[2][4] ));
   NOR2 \mult_19_2/AN1_2_3  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[2][3] ));
   NOR2 \mult_19_2/AN1_2_2  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[2][2] ));
   NOR2 \mult_19_2/AN1_2_1  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[2][1] ));
   NOR2 \mult_19_2/AN1_2_0_0  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[2][0] ));
   NOR2 \mult_19_2/AN2_1_7  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[1][7] ));
   NOR2 \mult_19_2/AN1_1_6  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[1][6] ));
   NOR2 \mult_19_2/AN1_1_5  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[1][5] ));
   NOR2 \mult_19_2/AN1_1_4  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[1][4] ));
   NOR2 \mult_19_2/AN1_1_3  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[1][3] ));
   NOR2 \mult_19_2/AN1_1_2  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[1][2] ));
   NOR2 \mult_19_2/AN1_1_1  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[1][1] ));
   NOR2 \mult_19_2/AN1_1_0_0  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[1][0] ));
   NOR2 \mult_19_2/AN2_0_7  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[0][7] ));
   NOR2 \mult_19_2/AN1_0_6  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[0][6] ));
   NOR2 \mult_19_2/AN1_0_5  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[0][5] ));
   NOR2 \mult_19_2/AN1_0_4  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[0][4] ));
   NOR2 \mult_19_2/AN1_0_3  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[0][3] ));
   NOR2 \mult_19_2/AN1_0_2  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[0][2] ));
   NOR2 \mult_19_2/AN1_0_1  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[0][1] ));
   NOR2 \mult_19_2/AN1_0_0_0  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(N17));
   OAI21 \mult_19/FS_1/U6_1_0_3  (.OUT(\mult_19/FS_1/C[1][3][0] ),
	.C(n2875),
	.B(n2874),
	.A(n2873));
   OAI21 \mult_19/FS_1/U6_0_3_1  (.OUT(\mult_19/FS_1/C[1][3][1] ),
	.C(\mult_19/FS_1/G_n_int[0][3][0] ),
	.B(n2871),
	.A(n2870));
   XOR2 \mult_19/FS_1/U3_C_0_3_1  (.A(\mult_19/FS_1/PG_int[0][3][1] ),
	.B(\mult_19/FS_1/C[1][3][1] ),
	.OUT(N16));
   XOR2 \mult_19/FS_1/U3_C_0_3_0  (.A(\mult_19/FS_1/PG_int[0][3][0] ),
	.B(\mult_19/FS_1/C[1][3][0] ),
	.OUT(N15));
   NAND2 \mult_19/FS_1/U3_B_0_3_0  (.A(\mult_19/FS_1/G_n_int[0][3][0] ),
	.B(\mult_19/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2867));
   NAND2 \mult_19/FS_1/U2_0_3_0  (.A(\mult_19/A1[12] ),
	.B(\mult_19/A2[12] ),
	.OUT(\mult_19/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_19/FS_1/U1_0_3_0  (.A(n2865),
	.B(n2866),
	.OUT(\mult_19/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_19/FS_1/U6_0_2_3  (.OUT(\mult_19/FS_1/C[1][2][3] ),
	.C(\mult_19/FS_1/G_n_int[0][2][2] ),
	.B(n2864),
	.A(n2863));
   OAI21 \mult_19/FS_1/U5_0_2_3  (.OUT(\mult_19/FS_1/G[1][0][2] ),
	.C(\mult_19/FS_1/G_n_int[0][2][3] ),
	.B(n2862),
	.A(n2861));
   NAND2 \mult_19/FS_1/U4_0_2_3  (.A(\mult_19/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_19/FS_1/P[0][2][3] ),
	.OUT(n2874));
   XOR2 \mult_19/FS_1/U3_C_0_2_3  (.A(\mult_19/FS_1/PG_int[0][2][3] ),
	.B(\mult_19/FS_1/C[1][2][3] ),
	.OUT(N14));
   NAND2 \mult_19/FS_1/U3_B_0_2_3  (.A(\mult_19/FS_1/G_n_int[0][2][3] ),
	.B(\mult_19/FS_1/P[0][2][3] ),
	.OUT(n2860));
   NAND2 \mult_19/FS_1/U2_0_2_3  (.A(\mult_19/A1[11] ),
	.B(\mult_19/A2[11] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_19/FS_1/U1_0_2_3  (.A(n2858),
	.B(n2859),
	.OUT(\mult_19/FS_1/P[0][2][3] ));
   OAI21 \mult_19/FS_1/U6_0_2_2  (.OUT(\mult_19/FS_1/C[1][2][2] ),
	.C(\mult_19/FS_1/G_n_int[0][2][1] ),
	.B(n2857),
	.A(n2856));
   OAI21 \mult_19/FS_1/U5_0_2_2  (.OUT(\mult_19/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_19/FS_1/G_n_int[0][2][2] ),
	.B(n2864),
	.A(n2855));
   NAND2 \mult_19/FS_1/U4_0_2_2  (.A(\mult_19/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_19/FS_1/P[0][2][2] ),
	.OUT(n2854));
   XOR2 \mult_19/FS_1/U3_C_0_2_2  (.A(\mult_19/FS_1/PG_int[0][2][2] ),
	.B(\mult_19/FS_1/C[1][2][2] ),
	.OUT(N13));
   NAND2 \mult_19/FS_1/U3_B_0_2_2  (.A(\mult_19/FS_1/G_n_int[0][2][2] ),
	.B(\mult_19/FS_1/P[0][2][2] ),
	.OUT(n2853));
   NAND2 \mult_19/FS_1/U2_0_2_2  (.A(\mult_19/A1[10] ),
	.B(\mult_19/A2[10] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_19/FS_1/U1_0_2_2  (.A(n2851),
	.B(n2852),
	.OUT(\mult_19/FS_1/P[0][2][2] ));
   OAI21 \mult_19/FS_1/U6_0_2_1  (.OUT(\mult_19/FS_1/C[1][2][1] ),
	.C(\mult_19/FS_1/G_n_int[0][2][0] ),
	.B(n2850),
	.A(n2873));
   OAI21 \mult_19/FS_1/U5_0_2_1  (.OUT(\mult_19/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_19/FS_1/G_n_int[0][2][1] ),
	.B(n2857),
	.A(\mult_19/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19/FS_1/U4_0_2_1  (.A(\mult_19/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_19/FS_1/P[0][2][1] ),
	.OUT(n2849));
   XOR2 \mult_19/FS_1/U3_C_0_2_1  (.A(\mult_19/FS_1/PG_int[0][2][1] ),
	.B(\mult_19/FS_1/C[1][2][1] ),
	.OUT(N12));
   NAND2 \mult_19/FS_1/U3_B_0_2_1  (.A(\mult_19/FS_1/G_n_int[0][2][1] ),
	.B(\mult_19/FS_1/P[0][2][1] ),
	.OUT(n2848));
   NAND2 \mult_19/FS_1/U2_0_2_1  (.A(\mult_19/A1[9] ),
	.B(\mult_19/A2[9] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_19/FS_1/U1_0_2_1  (.A(n2846),
	.B(n2847),
	.OUT(\mult_19/FS_1/P[0][2][1] ));
   XOR2 \mult_19/FS_1/U3_C_0_2_0  (.A(\mult_19/FS_1/PG_int[0][2][0] ),
	.B(\mult_19/FS_1/C[1][2][0] ),
	.OUT(N11));
   NAND2 \mult_19/FS_1/U3_B_0_2_0  (.A(\mult_19/FS_1/G_n_int[0][2][0] ),
	.B(\mult_19/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2845));
   NAND2 \mult_19/FS_1/U2_0_2_0  (.A(\mult_19/A1[8] ),
	.B(\mult_19/A2[8] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19/FS_1/U1_0_2_0  (.A(n2843),
	.B(n2844),
	.OUT(\mult_19/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_19/FS_1/U3_B_0_1_3  (.A(\mult_19/FS_1/G_n_int[0][1][3] ),
	.B(\mult_19/FS_1/P[0][1][3] ),
	.OUT(n2842));
   NAND2 \mult_19/FS_1/U2_0_1_3  (.A(\mult_19/A1[7] ),
	.B(\mult_19/A2[7] ),
	.OUT(\mult_19/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_19/FS_1/U1_0_1_3  (.A(n2840),
	.B(n2841),
	.OUT(\mult_19/FS_1/P[0][1][3] ));
   inverter \mult_19/AN1_7  (.IN(matrix00[7]),
	.OUT(\mult_19/A_not[7] ));
   inverter \mult_19/AN1_6  (.IN(matrix00[6]),
	.OUT(\mult_19/A_notx [6]));
   inverter \mult_19/AN1_5  (.IN(matrix00[5]),
	.OUT(\mult_19/A_notx [5]));
   inverter \mult_19/AN1_4  (.IN(matrix00[4]),
	.OUT(\mult_19/A_notx [4]));
   inverter \mult_19/AN1_3  (.IN(matrix00[3]),
	.OUT(\mult_19/A_notx [3]));
   inverter \mult_19/AN1_2  (.IN(matrix00[2]),
	.OUT(\mult_19/A_notx [2]));
   inverter \mult_19/AN1_1  (.IN(matrix00[1]),
	.OUT(\mult_19/A_notx [1]));
   inverter \mult_19/AN1_0  (.IN(matrix00[0]),
	.OUT(\mult_19/A_notx [0]));
   inverter \mult_19/AN1_7_0  (.IN(vector_0[7]),
	.OUT(\mult_19/B_not[7] ));
   inverter \mult_19/AN1_6_0  (.IN(vector_0[6]),
	.OUT(\mult_19/B_notx [6]));
   inverter \mult_19/AN1_5_0  (.IN(vector_0[5]),
	.OUT(\mult_19/B_notx [5]));
   inverter \mult_19/AN1_4_0  (.IN(vector_0[4]),
	.OUT(\mult_19/B_notx [4]));
   inverter \mult_19/AN1_3_0  (.IN(vector_0[3]),
	.OUT(\mult_19/B_notx [3]));
   inverter \mult_19/AN1_2_0  (.IN(vector_0[2]),
	.OUT(\mult_19/B_notx [2]));
   inverter \mult_19/AN1_1_0  (.IN(vector_0[1]),
	.OUT(\mult_19/B_notx [1]));
   inverter \mult_19/AN1_0_0  (.IN(vector_0[0]),
	.OUT(\mult_19/B_notx [0]));
   NOR2 \mult_19/AN1_7_7  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[7][7] ));
   NOR2 \mult_19/AN3_7_6  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[7][6] ));
   NOR2 \mult_19/AN3_7_5  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[7][5] ));
   NOR2 \mult_19/AN3_7_4  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[7][4] ));
   NOR2 \mult_19/AN3_7_3  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[7][3] ));
   NOR2 \mult_19/AN3_7_2  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[7][2] ));
   NOR2 \mult_19/AN3_7_1  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[7][1] ));
   NOR2 \mult_19/AN3_7_0  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[7][0] ));
   NOR2 \mult_19/AN2_6_7  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[6][7] ));
   NOR2 \mult_19/AN1_6_6  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[6][6] ));
   NOR2 \mult_19/AN1_6_5  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[6][5] ));
   NOR2 \mult_19/AN1_6_4  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[6][4] ));
   NOR2 \mult_19/AN1_6_3  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[6][3] ));
   NOR2 \mult_19/AN1_6_2  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[6][2] ));
   NOR2 \mult_19/AN1_6_1  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[6][1] ));
   NOR2 \mult_19/AN1_6_0_0  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[6][0] ));
   NOR2 \mult_19/AN2_5_7  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[5][7] ));
   NOR2 \mult_19/AN1_5_6  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[5][6] ));
   NOR2 \mult_19/AN1_5_5  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[5][5] ));
   NOR2 \mult_19/AN1_5_4  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[5][4] ));
   NOR2 \mult_19/AN1_5_3  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[5][3] ));
   NOR2 \mult_19/AN1_5_2  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[5][2] ));
   NOR2 \mult_19/AN1_5_1  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[5][1] ));
   NOR2 \mult_19/AN1_5_0_0  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[5][0] ));
   NOR2 \mult_19/AN2_4_7  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[4][7] ));
   NOR2 \mult_19/AN1_4_6  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[4][6] ));
   NOR2 \mult_19/AN1_4_5  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[4][5] ));
   NOR2 \mult_19/AN1_4_4  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[4][4] ));
   NOR2 \mult_19/AN1_4_3  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[4][3] ));
   NOR2 \mult_19/AN1_4_2  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[4][2] ));
   NOR2 \mult_19/AN1_4_1  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[4][1] ));
   NOR2 \mult_19/AN1_4_0_0  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[4][0] ));
   NOR2 \mult_19/AN2_3_7  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[3][7] ));
   NOR2 \mult_19/AN1_3_6  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[3][6] ));
   NOR2 \mult_19/AN1_3_5  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[3][5] ));
   NOR2 \mult_19/AN1_3_4  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[3][4] ));
   NOR2 \mult_19/AN1_3_3  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[3][3] ));
   NOR2 \mult_19/AN1_3_2  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[3][2] ));
   NOR2 \mult_19/AN1_3_1  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[3][1] ));
   NOR2 \mult_19/AN1_3_0_0  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[3][0] ));
   NOR2 \mult_19/AN2_2_7  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[2][7] ));
   NOR2 \mult_19/AN1_2_6  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[2][6] ));
   NOR2 \mult_19/AN1_2_5  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[2][5] ));
   NOR2 \mult_19/AN1_2_4  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[2][4] ));
   NOR2 \mult_19/AN1_2_3  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[2][3] ));
   NOR2 \mult_19/AN1_2_2  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[2][2] ));
   NOR2 \mult_19/AN1_2_1  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[2][1] ));
   NOR2 \mult_19/AN1_2_0_0  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[2][0] ));
   NOR2 \mult_19/AN2_1_7  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[1][7] ));
   NOR2 \mult_19/AN1_1_6  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[1][6] ));
   NOR2 \mult_19/AN1_1_5  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[1][5] ));
   NOR2 \mult_19/AN1_1_4  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[1][4] ));
   NOR2 \mult_19/AN1_1_3  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[1][3] ));
   NOR2 \mult_19/AN1_1_2  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[1][2] ));
   NOR2 \mult_19/AN1_1_1  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[1][1] ));
   NOR2 \mult_19/AN1_1_0_0  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[1][0] ));
   NOR2 \mult_19/AN2_0_7  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[0][7] ));
   NOR2 \mult_19/AN1_0_6  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[0][6] ));
   NOR2 \mult_19/AN1_0_5  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[0][5] ));
   NOR2 \mult_19/AN1_0_4  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[0][4] ));
   NOR2 \mult_19/AN1_0_3  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[0][3] ));
   NOR2 \mult_19/AN1_0_2  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[0][2] ));
   NOR2 \mult_19/AN1_0_1  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[0][1] ));
   NOR2 \mult_19/AN1_0_0_0  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [0]),
	.OUT(N1));
   inverter U19 (.IN(clk),
	.OUT(n17));
   inverter U20 (.IN(clk),
	.OUT(n18));
   inverter U21 (.IN(clk),
	.OUT(n19));
   inverter U22 (.IN(clk),
	.OUT(n20));
   inverter U23 (.IN(clk),
	.OUT(n21));
   inverter U24 (.IN(clk),
	.OUT(n22));
   inverter U25 (.IN(clk),
	.OUT(n23));
   inverter U26 (.IN(clk),
	.OUT(n24));
   inverter U27 (.IN(clk),
	.OUT(n25));
   inverter U28 (.IN(clk),
	.OUT(n26));
   inverter U29 (.IN(clk),
	.OUT(n27));
   inverter U30 (.IN(clk),
	.OUT(n28));
   inverter U31 (.IN(clk),
	.OUT(n29));
   inverter U32 (.IN(clk),
	.OUT(n30));
   inverter U33 (.IN(clk),
	.OUT(n31));
   inverter U34 (.IN(clk),
	.OUT(n32));
   inverter U35 (.IN(clk),
	.OUT(n33));
   inverter U36 (.IN(clk),
	.OUT(n34));
   inverter U37 (.IN(clk),
	.OUT(n35));
   inverter U38 (.IN(clk),
	.OUT(n36));
   inverter U39 (.IN(clk),
	.OUT(n37));
   inverter U40 (.IN(clk),
	.OUT(n38));
   inverter U41 (.IN(clk),
	.OUT(n39));
   inverter U42 (.IN(clk),
	.OUT(n40));
   inverter U43 (.IN(clk),
	.OUT(n41));
   inverter U44 (.IN(clk),
	.OUT(n42));
   inverter U45 (.IN(clk),
	.OUT(n43));
   inverter U46 (.IN(clk),
	.OUT(n44));
   inverter U47 (.IN(clk),
	.OUT(n45));
   inverter U48 (.IN(clk),
	.OUT(n46));
   inverter U49 (.IN(clk),
	.OUT(n47));
   inverter U50 (.IN(clk),
	.OUT(n48));
   inverter U51 (.IN(clk),
	.OUT(n49));
   inverter U52 (.IN(clk),
	.OUT(n50));
   inverter U53 (.IN(clk),
	.OUT(n51));
   inverter U54 (.IN(clk),
	.OUT(n52));
   inverter U55 (.IN(clk),
	.OUT(n53));
   inverter U56 (.IN(rst_n),
	.OUT(n54));
   inverter U57 (.IN(rst_n),
	.OUT(n55));
   inverter U58 (.IN(clk),
	.OUT(n56));
   inverter U59 (.IN(clk),
	.OUT(n57));
   inverter U60 (.IN(clk),
	.OUT(n58));
   inverter U61 (.IN(clk),
	.OUT(n59));
   inverter U62 (.IN(clk),
	.OUT(n60));
   inverter U63 (.IN(clk),
	.OUT(n61));
   inverter U64 (.IN(clk),
	.OUT(n62));
   inverter U65 (.IN(clk),
	.OUT(n63));
   inverter U66 (.IN(clk),
	.OUT(n64));
   inverter U67 (.IN(clk),
	.OUT(n65));
   inverter U68 (.IN(n2826),
	.OUT(\mult_19/FS_1/TEMP_P[0][0][0] ));
   inverter U69 (.IN(n2876),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][0][0] ));
   inverter U70 (.IN(n2926),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][0][0] ));
   inverter U71 (.IN(n2976),
	.OUT(\mult_20/FS_1/TEMP_P[0][0][0] ));
   inverter U72 (.IN(n3026),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][0][0] ));
   inverter U73 (.IN(n3076),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][0][0] ));
   inverter U74 (.IN(n3126),
	.OUT(\mult_21/FS_1/TEMP_P[0][0][0] ));
   inverter U75 (.IN(n3176),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][0][0] ));
   inverter U76 (.IN(n3226),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][0][0] ));
   inverter U77 (.IN(\mult_21_3/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3227));
   inverter U78 (.IN(n3228),
	.OUT(\mult_21_3/FS_1/P[0][0][1] ));
   inverter U79 (.IN(\mult_21_3/FS_1/P[0][0][1] ),
	.OUT(n3229));
   inverter U80 (.IN(n3230),
	.OUT(\mult_21_3/FS_1/P[0][0][2] ));
   inverter U81 (.IN(\mult_21_3/FS_1/P[0][0][2] ),
	.OUT(n3231));
   inverter U82 (.IN(n3232),
	.OUT(\mult_21_3/FS_1/P[0][0][3] ));
   inverter U83 (.IN(\mult_21_3/FS_1/P[0][0][3] ),
	.OUT(n3233));
   inverter U84 (.IN(n3272),
	.OUT(\mult_21_3/FS_1/C[1][2][0] ));
   inverter U85 (.IN(n3234),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][1][0] ));
   inverter U86 (.IN(\mult_21_3/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3235));
   inverter U87 (.IN(n3236),
	.OUT(\mult_21_3/FS_1/P[0][1][1] ));
   inverter U88 (.IN(n3268),
	.OUT(\mult_21_3/FS_1/P[0][3][1] ));
   inverter U89 (.IN(\mult_21_3/FS_1/P[0][3][1] ),
	.OUT(n3269));
   inverter U90 (.IN(\mult_21_3/FS_1/P[0][1][1] ),
	.OUT(n3237));
   inverter U91 (.IN(n3238),
	.OUT(\mult_21_3/FS_1/P[0][1][2] ));
   inverter U92 (.IN(\mult_21_3/FS_1/P[0][1][2] ),
	.OUT(n3239));
   inverter U93 (.IN(\mult_21_3/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_21_3/FS_1/G[1][0][1] ));
   inverter U94 (.IN(\mult_21_2/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3177));
   inverter U95 (.IN(n3178),
	.OUT(\mult_21_2/FS_1/P[0][0][1] ));
   inverter U96 (.IN(\mult_21_2/FS_1/P[0][0][1] ),
	.OUT(n3179));
   inverter U97 (.IN(n3180),
	.OUT(\mult_21_2/FS_1/P[0][0][2] ));
   inverter U98 (.IN(\mult_21_2/FS_1/P[0][0][2] ),
	.OUT(n3181));
   inverter U99 (.IN(n3182),
	.OUT(\mult_21_2/FS_1/P[0][0][3] ));
   inverter U100 (.IN(\mult_21_2/FS_1/P[0][0][3] ),
	.OUT(n3183));
   inverter U101 (.IN(n3222),
	.OUT(\mult_21_2/FS_1/C[1][2][0] ));
   inverter U102 (.IN(n3184),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][1][0] ));
   inverter U103 (.IN(\mult_21_2/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3185));
   inverter U104 (.IN(n3186),
	.OUT(\mult_21_2/FS_1/P[0][1][1] ));
   inverter U105 (.IN(n3218),
	.OUT(\mult_21_2/FS_1/P[0][3][1] ));
   inverter U106 (.IN(\mult_21_2/FS_1/P[0][3][1] ),
	.OUT(n3219));
   inverter U107 (.IN(\mult_21_2/FS_1/P[0][1][1] ),
	.OUT(n3187));
   inverter U108 (.IN(n3188),
	.OUT(\mult_21_2/FS_1/P[0][1][2] ));
   inverter U109 (.IN(\mult_21_2/FS_1/P[0][1][2] ),
	.OUT(n3189));
   inverter U110 (.IN(\mult_21_2/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_21_2/FS_1/G[1][0][1] ));
   inverter U111 (.IN(\mult_21/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3127));
   inverter U112 (.IN(n3128),
	.OUT(\mult_21/FS_1/P[0][0][1] ));
   inverter U113 (.IN(\mult_21/FS_1/P[0][0][1] ),
	.OUT(n3129));
   inverter U114 (.IN(n3130),
	.OUT(\mult_21/FS_1/P[0][0][2] ));
   inverter U115 (.IN(\mult_21/FS_1/P[0][0][2] ),
	.OUT(n3131));
   inverter U116 (.IN(n3132),
	.OUT(\mult_21/FS_1/P[0][0][3] ));
   inverter U117 (.IN(\mult_21/FS_1/P[0][0][3] ),
	.OUT(n3133));
   inverter U118 (.IN(n3172),
	.OUT(\mult_21/FS_1/C[1][2][0] ));
   inverter U119 (.IN(n3134),
	.OUT(\mult_21/FS_1/TEMP_P[0][1][0] ));
   inverter U120 (.IN(\mult_21/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3135));
   inverter U121 (.IN(n3136),
	.OUT(\mult_21/FS_1/P[0][1][1] ));
   inverter U122 (.IN(n3168),
	.OUT(\mult_21/FS_1/P[0][3][1] ));
   inverter U123 (.IN(\mult_21/FS_1/P[0][3][1] ),
	.OUT(n3169));
   inverter U124 (.IN(\mult_21/FS_1/P[0][1][1] ),
	.OUT(n3137));
   inverter U125 (.IN(n3138),
	.OUT(\mult_21/FS_1/P[0][1][2] ));
   inverter U126 (.IN(\mult_21/FS_1/P[0][1][2] ),
	.OUT(n3139));
   inverter U127 (.IN(\mult_21/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_21/FS_1/G[1][0][1] ));
   inverter U128 (.IN(\mult_20_3/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3077));
   inverter U129 (.IN(n3078),
	.OUT(\mult_20_3/FS_1/P[0][0][1] ));
   inverter U130 (.IN(\mult_20_3/FS_1/P[0][0][1] ),
	.OUT(n3079));
   inverter U131 (.IN(n3080),
	.OUT(\mult_20_3/FS_1/P[0][0][2] ));
   inverter U132 (.IN(\mult_20_3/FS_1/P[0][0][2] ),
	.OUT(n3081));
   inverter U133 (.IN(n3082),
	.OUT(\mult_20_3/FS_1/P[0][0][3] ));
   inverter U134 (.IN(\mult_20_3/FS_1/P[0][0][3] ),
	.OUT(n3083));
   inverter U135 (.IN(n3122),
	.OUT(\mult_20_3/FS_1/C[1][2][0] ));
   inverter U136 (.IN(n3084),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][1][0] ));
   inverter U137 (.IN(\mult_20_3/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3085));
   inverter U138 (.IN(n3086),
	.OUT(\mult_20_3/FS_1/P[0][1][1] ));
   inverter U139 (.IN(n3118),
	.OUT(\mult_20_3/FS_1/P[0][3][1] ));
   inverter U140 (.IN(\mult_20_3/FS_1/P[0][3][1] ),
	.OUT(n3119));
   inverter U141 (.IN(\mult_20_3/FS_1/P[0][1][1] ),
	.OUT(n3087));
   inverter U142 (.IN(n3088),
	.OUT(\mult_20_3/FS_1/P[0][1][2] ));
   inverter U143 (.IN(\mult_20_3/FS_1/P[0][1][2] ),
	.OUT(n3089));
   inverter U144 (.IN(\mult_20_3/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_20_3/FS_1/G[1][0][1] ));
   inverter U145 (.IN(\mult_20_2/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3027));
   inverter U146 (.IN(n3028),
	.OUT(\mult_20_2/FS_1/P[0][0][1] ));
   inverter U147 (.IN(\mult_20_2/FS_1/P[0][0][1] ),
	.OUT(n3029));
   inverter U148 (.IN(n3030),
	.OUT(\mult_20_2/FS_1/P[0][0][2] ));
   inverter U149 (.IN(\mult_20_2/FS_1/P[0][0][2] ),
	.OUT(n3031));
   inverter U150 (.IN(n3032),
	.OUT(\mult_20_2/FS_1/P[0][0][3] ));
   inverter U151 (.IN(\mult_20_2/FS_1/P[0][0][3] ),
	.OUT(n3033));
   inverter U152 (.IN(n3072),
	.OUT(\mult_20_2/FS_1/C[1][2][0] ));
   inverter U153 (.IN(n3034),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][1][0] ));
   inverter U154 (.IN(\mult_20_2/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3035));
   inverter U155 (.IN(n3036),
	.OUT(\mult_20_2/FS_1/P[0][1][1] ));
   inverter U156 (.IN(n3068),
	.OUT(\mult_20_2/FS_1/P[0][3][1] ));
   inverter U157 (.IN(\mult_20_2/FS_1/P[0][3][1] ),
	.OUT(n3069));
   inverter U158 (.IN(\mult_20_2/FS_1/P[0][1][1] ),
	.OUT(n3037));
   inverter U159 (.IN(n3038),
	.OUT(\mult_20_2/FS_1/P[0][1][2] ));
   inverter U160 (.IN(\mult_20_2/FS_1/P[0][1][2] ),
	.OUT(n3039));
   inverter U161 (.IN(\mult_20_2/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_20_2/FS_1/G[1][0][1] ));
   inverter U162 (.IN(\mult_20/FS_1/TEMP_P[0][0][0] ),
	.OUT(n2977));
   inverter U163 (.IN(n2978),
	.OUT(\mult_20/FS_1/P[0][0][1] ));
   inverter U164 (.IN(\mult_20/FS_1/P[0][0][1] ),
	.OUT(n2979));
   inverter U165 (.IN(n2980),
	.OUT(\mult_20/FS_1/P[0][0][2] ));
   inverter U166 (.IN(\mult_20/FS_1/P[0][0][2] ),
	.OUT(n2981));
   inverter U167 (.IN(n2982),
	.OUT(\mult_20/FS_1/P[0][0][3] ));
   inverter U168 (.IN(\mult_20/FS_1/P[0][0][3] ),
	.OUT(n2983));
   inverter U169 (.IN(n3022),
	.OUT(\mult_20/FS_1/C[1][2][0] ));
   inverter U170 (.IN(n2984),
	.OUT(\mult_20/FS_1/TEMP_P[0][1][0] ));
   inverter U171 (.IN(\mult_20/FS_1/TEMP_P[0][1][0] ),
	.OUT(n2985));
   inverter U172 (.IN(n2986),
	.OUT(\mult_20/FS_1/P[0][1][1] ));
   inverter U173 (.IN(n3018),
	.OUT(\mult_20/FS_1/P[0][3][1] ));
   inverter U174 (.IN(\mult_20/FS_1/P[0][3][1] ),
	.OUT(n3019));
   inverter U175 (.IN(\mult_20/FS_1/P[0][1][1] ),
	.OUT(n2987));
   inverter U176 (.IN(n2988),
	.OUT(\mult_20/FS_1/P[0][1][2] ));
   inverter U177 (.IN(\mult_20/FS_1/P[0][1][2] ),
	.OUT(n2989));
   inverter U178 (.IN(\mult_20/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_20/FS_1/G[1][0][1] ));
   inverter U179 (.IN(\mult_19_3/FS_1/TEMP_P[0][0][0] ),
	.OUT(n2927));
   inverter U180 (.IN(n2928),
	.OUT(\mult_19_3/FS_1/P[0][0][1] ));
   inverter U181 (.IN(\mult_19_3/FS_1/P[0][0][1] ),
	.OUT(n2929));
   inverter U182 (.IN(n2930),
	.OUT(\mult_19_3/FS_1/P[0][0][2] ));
   inverter U183 (.IN(\mult_19_3/FS_1/P[0][0][2] ),
	.OUT(n2931));
   inverter U184 (.IN(n2932),
	.OUT(\mult_19_3/FS_1/P[0][0][3] ));
   inverter U185 (.IN(\mult_19_3/FS_1/P[0][0][3] ),
	.OUT(n2933));
   inverter U186 (.IN(n2972),
	.OUT(\mult_19_3/FS_1/C[1][2][0] ));
   inverter U187 (.IN(n2934),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][1][0] ));
   inverter U188 (.IN(\mult_19_3/FS_1/TEMP_P[0][1][0] ),
	.OUT(n2935));
   inverter U189 (.IN(n2936),
	.OUT(\mult_19_3/FS_1/P[0][1][1] ));
   inverter U190 (.IN(n2968),
	.OUT(\mult_19_3/FS_1/P[0][3][1] ));
   inverter U191 (.IN(\mult_19_3/FS_1/P[0][3][1] ),
	.OUT(n2969));
   inverter U192 (.IN(\mult_19_3/FS_1/P[0][1][1] ),
	.OUT(n2937));
   inverter U193 (.IN(n2938),
	.OUT(\mult_19_3/FS_1/P[0][1][2] ));
   inverter U194 (.IN(\mult_19_3/FS_1/P[0][1][2] ),
	.OUT(n2939));
   inverter U195 (.IN(\mult_19_3/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_19_3/FS_1/G[1][0][1] ));
   inverter U196 (.IN(\mult_19_2/FS_1/TEMP_P[0][0][0] ),
	.OUT(n2877));
   inverter U197 (.IN(n2878),
	.OUT(\mult_19_2/FS_1/P[0][0][1] ));
   inverter U198 (.IN(\mult_19_2/FS_1/P[0][0][1] ),
	.OUT(n2879));
   inverter U199 (.IN(n2880),
	.OUT(\mult_19_2/FS_1/P[0][0][2] ));
   inverter U200 (.IN(\mult_19_2/FS_1/P[0][0][2] ),
	.OUT(n2881));
   inverter U201 (.IN(n2882),
	.OUT(\mult_19_2/FS_1/P[0][0][3] ));
   inverter U202 (.IN(\mult_19_2/FS_1/P[0][0][3] ),
	.OUT(n2883));
   inverter U203 (.IN(n2922),
	.OUT(\mult_19_2/FS_1/C[1][2][0] ));
   inverter U204 (.IN(n2884),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][1][0] ));
   inverter U205 (.IN(\mult_19_2/FS_1/TEMP_P[0][1][0] ),
	.OUT(n2885));
   inverter U206 (.IN(n2886),
	.OUT(\mult_19_2/FS_1/P[0][1][1] ));
   inverter U207 (.IN(n2918),
	.OUT(\mult_19_2/FS_1/P[0][3][1] ));
   inverter U208 (.IN(\mult_19_2/FS_1/P[0][3][1] ),
	.OUT(n2919));
   inverter U209 (.IN(\mult_19_2/FS_1/P[0][1][1] ),
	.OUT(n2887));
   inverter U210 (.IN(n2888),
	.OUT(\mult_19_2/FS_1/P[0][1][2] ));
   inverter U211 (.IN(\mult_19_2/FS_1/P[0][1][2] ),
	.OUT(n2889));
   inverter U212 (.IN(\mult_19_2/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_19_2/FS_1/G[1][0][1] ));
   inverter U213 (.IN(\mult_19/FS_1/TEMP_P[0][0][0] ),
	.OUT(n2827));
   inverter U214 (.IN(n2828),
	.OUT(\mult_19/FS_1/P[0][0][1] ));
   inverter U215 (.IN(\mult_19/FS_1/P[0][0][1] ),
	.OUT(n2829));
   inverter U216 (.IN(n2830),
	.OUT(\mult_19/FS_1/P[0][0][2] ));
   inverter U217 (.IN(\mult_19/FS_1/P[0][0][2] ),
	.OUT(n2831));
   inverter U218 (.IN(n2832),
	.OUT(\mult_19/FS_1/P[0][0][3] ));
   inverter U219 (.IN(\mult_19/FS_1/P[0][0][3] ),
	.OUT(n2833));
   inverter U220 (.IN(n2872),
	.OUT(\mult_19/FS_1/C[1][2][0] ));
   inverter U221 (.IN(n2834),
	.OUT(\mult_19/FS_1/TEMP_P[0][1][0] ));
   inverter U222 (.IN(\mult_19/FS_1/TEMP_P[0][1][0] ),
	.OUT(n2835));
   inverter U223 (.IN(n2836),
	.OUT(\mult_19/FS_1/P[0][1][1] ));
   inverter U224 (.IN(n2868),
	.OUT(\mult_19/FS_1/P[0][3][1] ));
   inverter U225 (.IN(\mult_19/FS_1/P[0][3][1] ),
	.OUT(n2869));
   inverter U226 (.IN(\mult_19/FS_1/P[0][1][1] ),
	.OUT(n2837));
   inverter U227 (.IN(n2838),
	.OUT(\mult_19/FS_1/P[0][1][2] ));
   inverter U228 (.IN(\mult_19/FS_1/P[0][1][2] ),
	.OUT(n2839));
   inverter U229 (.IN(\mult_19/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_19/FS_1/G[1][0][1] ));
   NOR2 U230 (.A(n66),
	.B(n67),
	.OUT(\mult_19/A2[13] ));
   NOR2 U231 (.A(n68),
	.B(n69),
	.OUT(\mult_19/A2[12] ));
   NAND2 U232 (.A(n71),
	.B(n72),
	.OUT(n70));
   NOR2 U233 (.A(n73),
	.B(n74),
	.OUT(\mult_19/A2[10] ));
   NOR2 U234 (.A(n75),
	.B(n76),
	.OUT(\mult_19/A2[9] ));
   NOR2 U235 (.A(n77),
	.B(n78),
	.OUT(\mult_19/A2[8] ));
   NOR2 U236 (.A(n79),
	.B(n80),
	.OUT(\mult_19/A2[7] ));
   NOR2 U237 (.A(n81),
	.B(n82),
	.OUT(\mult_19_2/A2[13] ));
   NOR2 U238 (.A(n83),
	.B(n84),
	.OUT(\mult_19_2/A2[12] ));
   NAND2 U239 (.A(n86),
	.B(n87),
	.OUT(n85));
   NOR2 U240 (.A(n88),
	.B(n89),
	.OUT(\mult_19_2/A2[10] ));
   NOR2 U241 (.A(n90),
	.B(n91),
	.OUT(\mult_19_2/A2[9] ));
   NOR2 U242 (.A(n92),
	.B(n93),
	.OUT(\mult_19_2/A2[8] ));
   NOR2 U243 (.A(n94),
	.B(n95),
	.OUT(\mult_19_2/A2[7] ));
   NOR2 U244 (.A(n96),
	.B(n97),
	.OUT(\mult_19_3/A2[13] ));
   NOR2 U245 (.A(n98),
	.B(n99),
	.OUT(\mult_19_3/A2[12] ));
   NAND2 U246 (.A(n101),
	.B(n102),
	.OUT(n100));
   NOR2 U247 (.A(n103),
	.B(n104),
	.OUT(\mult_19_3/A2[10] ));
   NOR2 U248 (.A(n105),
	.B(n106),
	.OUT(\mult_19_3/A2[9] ));
   NOR2 U249 (.A(n107),
	.B(n108),
	.OUT(\mult_19_3/A2[8] ));
   NOR2 U250 (.A(n109),
	.B(n110),
	.OUT(\mult_19_3/A2[7] ));
   NOR2 U251 (.A(n111),
	.B(n112),
	.OUT(\mult_20/A2[13] ));
   NOR2 U252 (.A(n113),
	.B(n114),
	.OUT(\mult_20/A2[12] ));
   NAND2 U253 (.A(n116),
	.B(n117),
	.OUT(n115));
   NOR2 U254 (.A(n118),
	.B(n119),
	.OUT(\mult_20/A2[10] ));
   NOR2 U255 (.A(n120),
	.B(n121),
	.OUT(\mult_20/A2[9] ));
   NOR2 U256 (.A(n122),
	.B(n123),
	.OUT(\mult_20/A2[8] ));
   NOR2 U257 (.A(n124),
	.B(n125),
	.OUT(\mult_20/A2[7] ));
   NOR2 U258 (.A(n126),
	.B(n127),
	.OUT(\mult_20_2/A2[13] ));
   NOR2 U259 (.A(n128),
	.B(n129),
	.OUT(\mult_20_2/A2[12] ));
   NAND2 U260 (.A(n131),
	.B(n132),
	.OUT(n130));
   NOR2 U261 (.A(n133),
	.B(n134),
	.OUT(\mult_20_2/A2[10] ));
   NOR2 U262 (.A(n135),
	.B(n136),
	.OUT(\mult_20_2/A2[9] ));
   NOR2 U263 (.A(n137),
	.B(n138),
	.OUT(\mult_20_2/A2[8] ));
   NOR2 U264 (.A(n139),
	.B(n140),
	.OUT(\mult_20_2/A2[7] ));
   NOR2 U265 (.A(n141),
	.B(n142),
	.OUT(\mult_20_3/A2[13] ));
   NOR2 U266 (.A(n143),
	.B(n144),
	.OUT(\mult_20_3/A2[12] ));
   NAND2 U267 (.A(n146),
	.B(n147),
	.OUT(n145));
   NOR2 U268 (.A(n148),
	.B(n149),
	.OUT(\mult_20_3/A2[10] ));
   NOR2 U269 (.A(n150),
	.B(n151),
	.OUT(\mult_20_3/A2[9] ));
   NOR2 U270 (.A(n152),
	.B(n153),
	.OUT(\mult_20_3/A2[8] ));
   NOR2 U271 (.A(n154),
	.B(n155),
	.OUT(\mult_20_3/A2[7] ));
   NOR2 U272 (.A(n156),
	.B(n157),
	.OUT(\mult_21/A2[13] ));
   NOR2 U273 (.A(n158),
	.B(n159),
	.OUT(\mult_21/A2[12] ));
   NAND2 U274 (.A(n161),
	.B(n162),
	.OUT(n160));
   NOR2 U275 (.A(n163),
	.B(n164),
	.OUT(\mult_21/A2[10] ));
   NOR2 U276 (.A(n165),
	.B(n166),
	.OUT(\mult_21/A2[9] ));
   NOR2 U277 (.A(n167),
	.B(n168),
	.OUT(\mult_21/A2[8] ));
   NOR2 U278 (.A(n169),
	.B(n170),
	.OUT(\mult_21/A2[7] ));
   NOR2 U279 (.A(n171),
	.B(n172),
	.OUT(\mult_21_2/A2[13] ));
   NOR2 U280 (.A(n173),
	.B(n174),
	.OUT(\mult_21_2/A2[12] ));
   NAND2 U281 (.A(n176),
	.B(n177),
	.OUT(n175));
   NOR2 U282 (.A(n178),
	.B(n179),
	.OUT(\mult_21_2/A2[10] ));
   NOR2 U283 (.A(n180),
	.B(n181),
	.OUT(\mult_21_2/A2[9] ));
   NOR2 U284 (.A(n182),
	.B(n183),
	.OUT(\mult_21_2/A2[8] ));
   NOR2 U285 (.A(n184),
	.B(n185),
	.OUT(\mult_21_2/A2[7] ));
   NOR2 U286 (.A(n186),
	.B(n187),
	.OUT(\mult_21_3/A2[13] ));
   NOR2 U287 (.A(n188),
	.B(n189),
	.OUT(\mult_21_3/A2[12] ));
   NAND2 U288 (.A(n191),
	.B(n192),
	.OUT(n190));
   NOR2 U289 (.A(n193),
	.B(n194),
	.OUT(\mult_21_3/A2[10] ));
   NOR2 U290 (.A(n195),
	.B(n196),
	.OUT(\mult_21_3/A2[9] ));
   NOR2 U291 (.A(n197),
	.B(n198),
	.OUT(\mult_21_3/A2[8] ));
   NOR2 U292 (.A(n199),
	.B(n200),
	.OUT(\mult_21_3/A2[7] ));
   OAI21 U293 (.OUT(n201),
	.C(n202),
	.B(N31),
	.A(N15));
   AOI21 U294 (.OUT(n203),
	.C(n204),
	.B(N31),
	.A(N15));
   AOI21 U295 (.OUT(n205),
	.C(n208),
	.B(n207),
	.A(n206));
   AOI21 U296 (.OUT(n209),
	.C(n205),
	.B(n210),
	.A(N63));
   OAI21 U297 (.OUT(n211),
	.C(n212),
	.B(N191),
	.A(N175));
   AOI21 U298 (.OUT(n213),
	.C(n214),
	.B(N191),
	.A(N175));
   AOI21 U299 (.OUT(n215),
	.C(n218),
	.B(n217),
	.A(n216));
   AOI21 U300 (.OUT(n219),
	.C(n215),
	.B(n220),
	.A(N223));
   OAI21 U301 (.OUT(n221),
	.C(n222),
	.B(N111),
	.A(N95));
   AOI21 U302 (.OUT(n223),
	.C(n224),
	.B(N111),
	.A(N95));
   AOI21 U303 (.OUT(n225),
	.C(n228),
	.B(n227),
	.A(n226));
   AOI21 U304 (.OUT(n229),
	.C(n225),
	.B(n230),
	.A(N143));
   XOR2 U305 (.A(\mult_21_3/ab[1][7] ),
	.B(n232),
	.OUT(n231));
   XOR2 U306 (.A(\mult_21_3/ab[1][6] ),
	.B(\mult_21_3/ab[0][7] ),
	.OUT(n233));
   XOR2 U307 (.A(\mult_21_3/ab[1][5] ),
	.B(\mult_21_3/ab[0][6] ),
	.OUT(n234));
   XOR2 U308 (.A(n236),
	.B(n233),
	.OUT(n235));
   XOR2 U309 (.A(n238),
	.B(n239),
	.OUT(n237));
   XOR2 U310 (.A(\mult_21_3/ab[1][4] ),
	.B(\mult_21_3/ab[0][5] ),
	.OUT(n240));
   XOR2 U311 (.A(n242),
	.B(n234),
	.OUT(n241));
   XOR2 U312 (.A(\mult_21_3/ab[1][3] ),
	.B(\mult_21_3/ab[0][4] ),
	.OUT(n243));
   XOR2 U313 (.A(n245),
	.B(n240),
	.OUT(n244));
   XOR2 U314 (.A(n247),
	.B(n248),
	.OUT(n246));
   XOR2 U315 (.A(n250),
	.B(n251),
	.OUT(n249));
   XOR2 U316 (.A(n253),
	.B(n254),
	.OUT(n252));
   XOR2 U317 (.A(n256),
	.B(n257),
	.OUT(n255));
   XOR2 U318 (.A(n258),
	.B(n259),
	.OUT(n196));
   XOR2 U319 (.A(\mult_21_3/ab[1][2] ),
	.B(\mult_21_3/ab[0][3] ),
	.OUT(n260));
   XOR2 U320 (.A(n262),
	.B(n243),
	.OUT(n261));
   XOR2 U321 (.A(n264),
	.B(n265),
	.OUT(n263));
   XOR2 U322 (.A(n267),
	.B(n268),
	.OUT(n266));
   XOR2 U323 (.A(\mult_21_3/ab[1][1] ),
	.B(\mult_21_3/ab[0][2] ),
	.OUT(n269));
   XOR2 U324 (.A(n271),
	.B(n260),
	.OUT(n270));
   XOR2 U325 (.A(n273),
	.B(n274),
	.OUT(n272));
   XOR2 U326 (.A(n276),
	.B(n277),
	.OUT(n275));
   XOR2 U327 (.A(n279),
	.B(n280),
	.OUT(n278));
   XOR2 U328 (.A(n281),
	.B(n282),
	.OUT(n192));
   XOR2 U329 (.A(n195),
	.B(n196),
	.OUT(\mult_21_3/A1[8] ));
   XOR2 U330 (.A(n275),
	.B(n283),
	.OUT(\mult_21_3/A1[5] ));
   XOR2 U331 (.A(n272),
	.B(n284),
	.OUT(\mult_21_3/A1[3] ));
   XOR2 U332 (.A(n270),
	.B(n285),
	.OUT(\mult_21_3/A1[1] ));
   XOR2 U333 (.A(n187),
	.B(n186),
	.OUT(\mult_21_3/A1[12] ));
   XOR2 U334 (.A(n191),
	.B(n192),
	.OUT(\mult_21_3/A1[10] ));
   XOR2 U335 (.A(\mult_21_2/ab[1][7] ),
	.B(n287),
	.OUT(n286));
   XOR2 U336 (.A(\mult_21_2/ab[1][6] ),
	.B(\mult_21_2/ab[0][7] ),
	.OUT(n288));
   XOR2 U337 (.A(\mult_21_2/ab[1][5] ),
	.B(\mult_21_2/ab[0][6] ),
	.OUT(n289));
   XOR2 U338 (.A(n291),
	.B(n288),
	.OUT(n290));
   XOR2 U339 (.A(n293),
	.B(n294),
	.OUT(n292));
   XOR2 U340 (.A(\mult_21_2/ab[1][4] ),
	.B(\mult_21_2/ab[0][5] ),
	.OUT(n295));
   XOR2 U341 (.A(n297),
	.B(n289),
	.OUT(n296));
   XOR2 U342 (.A(\mult_21_2/ab[1][3] ),
	.B(\mult_21_2/ab[0][4] ),
	.OUT(n298));
   XOR2 U343 (.A(n300),
	.B(n295),
	.OUT(n299));
   XOR2 U344 (.A(n302),
	.B(n303),
	.OUT(n301));
   XOR2 U345 (.A(n305),
	.B(n306),
	.OUT(n304));
   XOR2 U346 (.A(n308),
	.B(n309),
	.OUT(n307));
   XOR2 U347 (.A(n311),
	.B(n312),
	.OUT(n310));
   XOR2 U348 (.A(n313),
	.B(n314),
	.OUT(n181));
   XOR2 U349 (.A(\mult_21_2/ab[1][2] ),
	.B(\mult_21_2/ab[0][3] ),
	.OUT(n315));
   XOR2 U350 (.A(n317),
	.B(n298),
	.OUT(n316));
   XOR2 U351 (.A(n319),
	.B(n320),
	.OUT(n318));
   XOR2 U352 (.A(n322),
	.B(n323),
	.OUT(n321));
   XOR2 U353 (.A(\mult_21_2/ab[1][1] ),
	.B(\mult_21_2/ab[0][2] ),
	.OUT(n324));
   XOR2 U354 (.A(n326),
	.B(n315),
	.OUT(n325));
   XOR2 U355 (.A(n328),
	.B(n329),
	.OUT(n327));
   XOR2 U356 (.A(n331),
	.B(n332),
	.OUT(n330));
   XOR2 U357 (.A(n334),
	.B(n335),
	.OUT(n333));
   XOR2 U358 (.A(n336),
	.B(n337),
	.OUT(n177));
   XOR2 U359 (.A(n180),
	.B(n181),
	.OUT(\mult_21_2/A1[8] ));
   XOR2 U360 (.A(n330),
	.B(n338),
	.OUT(\mult_21_2/A1[5] ));
   XOR2 U361 (.A(n327),
	.B(n339),
	.OUT(\mult_21_2/A1[3] ));
   XOR2 U362 (.A(n325),
	.B(n340),
	.OUT(\mult_21_2/A1[1] ));
   XOR2 U363 (.A(n172),
	.B(n171),
	.OUT(\mult_21_2/A1[12] ));
   XOR2 U364 (.A(n176),
	.B(n177),
	.OUT(\mult_21_2/A1[10] ));
   XOR2 U365 (.A(\mult_21/ab[1][7] ),
	.B(n342),
	.OUT(n341));
   XOR2 U366 (.A(\mult_21/ab[1][6] ),
	.B(\mult_21/ab[0][7] ),
	.OUT(n343));
   XOR2 U367 (.A(\mult_21/ab[1][5] ),
	.B(\mult_21/ab[0][6] ),
	.OUT(n344));
   XOR2 U368 (.A(n346),
	.B(n343),
	.OUT(n345));
   XOR2 U369 (.A(n348),
	.B(n349),
	.OUT(n347));
   XOR2 U370 (.A(\mult_21/ab[1][4] ),
	.B(\mult_21/ab[0][5] ),
	.OUT(n350));
   XOR2 U371 (.A(n352),
	.B(n344),
	.OUT(n351));
   XOR2 U372 (.A(\mult_21/ab[1][3] ),
	.B(\mult_21/ab[0][4] ),
	.OUT(n353));
   XOR2 U373 (.A(n355),
	.B(n350),
	.OUT(n354));
   XOR2 U374 (.A(n357),
	.B(n358),
	.OUT(n356));
   XOR2 U375 (.A(n360),
	.B(n361),
	.OUT(n359));
   XOR2 U376 (.A(n363),
	.B(n364),
	.OUT(n362));
   XOR2 U377 (.A(n366),
	.B(n367),
	.OUT(n365));
   XOR2 U378 (.A(n368),
	.B(n369),
	.OUT(n166));
   XOR2 U379 (.A(\mult_21/ab[1][2] ),
	.B(\mult_21/ab[0][3] ),
	.OUT(n370));
   XOR2 U380 (.A(n372),
	.B(n353),
	.OUT(n371));
   XOR2 U381 (.A(n374),
	.B(n375),
	.OUT(n373));
   XOR2 U382 (.A(n377),
	.B(n378),
	.OUT(n376));
   XOR2 U383 (.A(\mult_21/ab[1][1] ),
	.B(\mult_21/ab[0][2] ),
	.OUT(n379));
   XOR2 U384 (.A(n381),
	.B(n370),
	.OUT(n380));
   XOR2 U385 (.A(n383),
	.B(n384),
	.OUT(n382));
   XOR2 U386 (.A(n386),
	.B(n387),
	.OUT(n385));
   XOR2 U387 (.A(n389),
	.B(n390),
	.OUT(n388));
   XOR2 U388 (.A(n391),
	.B(n392),
	.OUT(n162));
   XOR2 U389 (.A(n165),
	.B(n166),
	.OUT(\mult_21/A1[8] ));
   XOR2 U390 (.A(n385),
	.B(n393),
	.OUT(\mult_21/A1[5] ));
   XOR2 U391 (.A(n382),
	.B(n394),
	.OUT(\mult_21/A1[3] ));
   XOR2 U392 (.A(n380),
	.B(n395),
	.OUT(\mult_21/A1[1] ));
   XOR2 U393 (.A(n157),
	.B(n156),
	.OUT(\mult_21/A1[12] ));
   XOR2 U394 (.A(n161),
	.B(n162),
	.OUT(\mult_21/A1[10] ));
   XOR2 U395 (.A(\mult_20_3/ab[1][7] ),
	.B(n397),
	.OUT(n396));
   XOR2 U396 (.A(\mult_20_3/ab[1][6] ),
	.B(\mult_20_3/ab[0][7] ),
	.OUT(n398));
   XOR2 U397 (.A(\mult_20_3/ab[1][5] ),
	.B(\mult_20_3/ab[0][6] ),
	.OUT(n399));
   XOR2 U398 (.A(n401),
	.B(n398),
	.OUT(n400));
   XOR2 U399 (.A(n403),
	.B(n404),
	.OUT(n402));
   XOR2 U400 (.A(\mult_20_3/ab[1][4] ),
	.B(\mult_20_3/ab[0][5] ),
	.OUT(n405));
   XOR2 U401 (.A(n407),
	.B(n399),
	.OUT(n406));
   XOR2 U402 (.A(\mult_20_3/ab[1][3] ),
	.B(\mult_20_3/ab[0][4] ),
	.OUT(n408));
   XOR2 U403 (.A(n410),
	.B(n405),
	.OUT(n409));
   XOR2 U404 (.A(n412),
	.B(n413),
	.OUT(n411));
   XOR2 U405 (.A(n415),
	.B(n416),
	.OUT(n414));
   XOR2 U406 (.A(n418),
	.B(n419),
	.OUT(n417));
   XOR2 U407 (.A(n421),
	.B(n422),
	.OUT(n420));
   XOR2 U408 (.A(n423),
	.B(n424),
	.OUT(n151));
   XOR2 U409 (.A(\mult_20_3/ab[1][2] ),
	.B(\mult_20_3/ab[0][3] ),
	.OUT(n425));
   XOR2 U410 (.A(n427),
	.B(n408),
	.OUT(n426));
   XOR2 U411 (.A(n429),
	.B(n430),
	.OUT(n428));
   XOR2 U412 (.A(n432),
	.B(n433),
	.OUT(n431));
   XOR2 U413 (.A(\mult_20_3/ab[1][1] ),
	.B(\mult_20_3/ab[0][2] ),
	.OUT(n434));
   XOR2 U414 (.A(n436),
	.B(n425),
	.OUT(n435));
   XOR2 U415 (.A(n438),
	.B(n439),
	.OUT(n437));
   XOR2 U416 (.A(n441),
	.B(n442),
	.OUT(n440));
   XOR2 U417 (.A(n444),
	.B(n445),
	.OUT(n443));
   XOR2 U418 (.A(n446),
	.B(n447),
	.OUT(n147));
   XOR2 U419 (.A(n150),
	.B(n151),
	.OUT(\mult_20_3/A1[8] ));
   XOR2 U420 (.A(n440),
	.B(n448),
	.OUT(\mult_20_3/A1[5] ));
   XOR2 U421 (.A(n437),
	.B(n449),
	.OUT(\mult_20_3/A1[3] ));
   XOR2 U422 (.A(n435),
	.B(n450),
	.OUT(\mult_20_3/A1[1] ));
   XOR2 U423 (.A(n142),
	.B(n141),
	.OUT(\mult_20_3/A1[12] ));
   XOR2 U424 (.A(n146),
	.B(n147),
	.OUT(\mult_20_3/A1[10] ));
   XOR2 U425 (.A(\mult_20_2/ab[1][7] ),
	.B(n452),
	.OUT(n451));
   XOR2 U426 (.A(\mult_20_2/ab[1][6] ),
	.B(\mult_20_2/ab[0][7] ),
	.OUT(n453));
   XOR2 U427 (.A(\mult_20_2/ab[1][5] ),
	.B(\mult_20_2/ab[0][6] ),
	.OUT(n454));
   XOR2 U428 (.A(n456),
	.B(n453),
	.OUT(n455));
   XOR2 U429 (.A(n458),
	.B(n459),
	.OUT(n457));
   XOR2 U430 (.A(\mult_20_2/ab[1][4] ),
	.B(\mult_20_2/ab[0][5] ),
	.OUT(n460));
   XOR2 U431 (.A(n462),
	.B(n454),
	.OUT(n461));
   XOR2 U432 (.A(\mult_20_2/ab[1][3] ),
	.B(\mult_20_2/ab[0][4] ),
	.OUT(n463));
   XOR2 U433 (.A(n465),
	.B(n460),
	.OUT(n464));
   XOR2 U434 (.A(n467),
	.B(n468),
	.OUT(n466));
   XOR2 U435 (.A(n470),
	.B(n471),
	.OUT(n469));
   XOR2 U436 (.A(n473),
	.B(n474),
	.OUT(n472));
   XOR2 U437 (.A(n476),
	.B(n477),
	.OUT(n475));
   XOR2 U438 (.A(n478),
	.B(n479),
	.OUT(n136));
   XOR2 U439 (.A(\mult_20_2/ab[1][2] ),
	.B(\mult_20_2/ab[0][3] ),
	.OUT(n480));
   XOR2 U440 (.A(n482),
	.B(n463),
	.OUT(n481));
   XOR2 U441 (.A(n484),
	.B(n485),
	.OUT(n483));
   XOR2 U442 (.A(n487),
	.B(n488),
	.OUT(n486));
   XOR2 U443 (.A(\mult_20_2/ab[1][1] ),
	.B(\mult_20_2/ab[0][2] ),
	.OUT(n489));
   XOR2 U444 (.A(n491),
	.B(n480),
	.OUT(n490));
   XOR2 U445 (.A(n493),
	.B(n494),
	.OUT(n492));
   XOR2 U446 (.A(n496),
	.B(n497),
	.OUT(n495));
   XOR2 U447 (.A(n499),
	.B(n500),
	.OUT(n498));
   XOR2 U448 (.A(n501),
	.B(n502),
	.OUT(n132));
   XOR2 U449 (.A(n135),
	.B(n136),
	.OUT(\mult_20_2/A1[8] ));
   XOR2 U450 (.A(n495),
	.B(n503),
	.OUT(\mult_20_2/A1[5] ));
   XOR2 U451 (.A(n492),
	.B(n504),
	.OUT(\mult_20_2/A1[3] ));
   XOR2 U452 (.A(n490),
	.B(n505),
	.OUT(\mult_20_2/A1[1] ));
   XOR2 U453 (.A(n127),
	.B(n126),
	.OUT(\mult_20_2/A1[12] ));
   XOR2 U454 (.A(n131),
	.B(n132),
	.OUT(\mult_20_2/A1[10] ));
   XOR2 U455 (.A(\mult_20/ab[1][7] ),
	.B(n507),
	.OUT(n506));
   XOR2 U456 (.A(\mult_20/ab[1][6] ),
	.B(\mult_20/ab[0][7] ),
	.OUT(n508));
   XOR2 U457 (.A(\mult_20/ab[1][5] ),
	.B(\mult_20/ab[0][6] ),
	.OUT(n509));
   XOR2 U458 (.A(n511),
	.B(n508),
	.OUT(n510));
   XOR2 U459 (.A(n513),
	.B(n514),
	.OUT(n512));
   XOR2 U460 (.A(\mult_20/ab[1][4] ),
	.B(\mult_20/ab[0][5] ),
	.OUT(n515));
   XOR2 U461 (.A(n517),
	.B(n509),
	.OUT(n516));
   XOR2 U462 (.A(\mult_20/ab[1][3] ),
	.B(\mult_20/ab[0][4] ),
	.OUT(n518));
   XOR2 U463 (.A(n520),
	.B(n515),
	.OUT(n519));
   XOR2 U464 (.A(n522),
	.B(n523),
	.OUT(n521));
   XOR2 U465 (.A(n525),
	.B(n526),
	.OUT(n524));
   XOR2 U466 (.A(n528),
	.B(n529),
	.OUT(n527));
   XOR2 U467 (.A(n531),
	.B(n532),
	.OUT(n530));
   XOR2 U468 (.A(n533),
	.B(n534),
	.OUT(n121));
   XOR2 U469 (.A(\mult_20/ab[1][2] ),
	.B(\mult_20/ab[0][3] ),
	.OUT(n535));
   XOR2 U470 (.A(n537),
	.B(n518),
	.OUT(n536));
   XOR2 U471 (.A(n539),
	.B(n540),
	.OUT(n538));
   XOR2 U472 (.A(n542),
	.B(n543),
	.OUT(n541));
   XOR2 U473 (.A(\mult_20/ab[1][1] ),
	.B(\mult_20/ab[0][2] ),
	.OUT(n544));
   XOR2 U474 (.A(n546),
	.B(n535),
	.OUT(n545));
   XOR2 U475 (.A(n548),
	.B(n549),
	.OUT(n547));
   XOR2 U476 (.A(n551),
	.B(n552),
	.OUT(n550));
   XOR2 U477 (.A(n554),
	.B(n555),
	.OUT(n553));
   XOR2 U478 (.A(n556),
	.B(n557),
	.OUT(n117));
   XOR2 U479 (.A(n120),
	.B(n121),
	.OUT(\mult_20/A1[8] ));
   XOR2 U480 (.A(n550),
	.B(n558),
	.OUT(\mult_20/A1[5] ));
   XOR2 U481 (.A(n547),
	.B(n559),
	.OUT(\mult_20/A1[3] ));
   XOR2 U482 (.A(n545),
	.B(n560),
	.OUT(\mult_20/A1[1] ));
   XOR2 U483 (.A(n112),
	.B(n111),
	.OUT(\mult_20/A1[12] ));
   XOR2 U484 (.A(n116),
	.B(n117),
	.OUT(\mult_20/A1[10] ));
   XOR2 U485 (.A(\mult_19_3/ab[1][7] ),
	.B(n562),
	.OUT(n561));
   XOR2 U486 (.A(\mult_19_3/ab[1][6] ),
	.B(\mult_19_3/ab[0][7] ),
	.OUT(n563));
   XOR2 U487 (.A(\mult_19_3/ab[1][5] ),
	.B(\mult_19_3/ab[0][6] ),
	.OUT(n564));
   XOR2 U488 (.A(n566),
	.B(n563),
	.OUT(n565));
   XOR2 U489 (.A(n568),
	.B(n569),
	.OUT(n567));
   XOR2 U490 (.A(\mult_19_3/ab[1][4] ),
	.B(\mult_19_3/ab[0][5] ),
	.OUT(n570));
   XOR2 U491 (.A(n572),
	.B(n564),
	.OUT(n571));
   XOR2 U492 (.A(\mult_19_3/ab[1][3] ),
	.B(\mult_19_3/ab[0][4] ),
	.OUT(n573));
   XOR2 U493 (.A(n575),
	.B(n570),
	.OUT(n574));
   XOR2 U494 (.A(n577),
	.B(n578),
	.OUT(n576));
   XOR2 U495 (.A(n580),
	.B(n581),
	.OUT(n579));
   XOR2 U496 (.A(n583),
	.B(n584),
	.OUT(n582));
   XOR2 U497 (.A(n586),
	.B(n587),
	.OUT(n585));
   XOR2 U498 (.A(n588),
	.B(n589),
	.OUT(n106));
   XOR2 U499 (.A(\mult_19_3/ab[1][2] ),
	.B(\mult_19_3/ab[0][3] ),
	.OUT(n590));
   XOR2 U500 (.A(n592),
	.B(n573),
	.OUT(n591));
   XOR2 U501 (.A(n594),
	.B(n595),
	.OUT(n593));
   XOR2 U502 (.A(n597),
	.B(n598),
	.OUT(n596));
   XOR2 U503 (.A(\mult_19_3/ab[1][1] ),
	.B(\mult_19_3/ab[0][2] ),
	.OUT(n599));
   XOR2 U504 (.A(n601),
	.B(n590),
	.OUT(n600));
   XOR2 U505 (.A(n603),
	.B(n604),
	.OUT(n602));
   XOR2 U506 (.A(n606),
	.B(n607),
	.OUT(n605));
   XOR2 U507 (.A(n609),
	.B(n610),
	.OUT(n608));
   XOR2 U508 (.A(n611),
	.B(n612),
	.OUT(n102));
   XOR2 U509 (.A(n105),
	.B(n106),
	.OUT(\mult_19_3/A1[8] ));
   XOR2 U510 (.A(n605),
	.B(n613),
	.OUT(\mult_19_3/A1[5] ));
   XOR2 U511 (.A(n602),
	.B(n614),
	.OUT(\mult_19_3/A1[3] ));
   XOR2 U512 (.A(n600),
	.B(n615),
	.OUT(\mult_19_3/A1[1] ));
   XOR2 U513 (.A(n97),
	.B(n96),
	.OUT(\mult_19_3/A1[12] ));
   XOR2 U514 (.A(n101),
	.B(n102),
	.OUT(\mult_19_3/A1[10] ));
   XOR2 U515 (.A(\mult_19_2/ab[1][7] ),
	.B(n617),
	.OUT(n616));
   XOR2 U516 (.A(\mult_19_2/ab[1][6] ),
	.B(\mult_19_2/ab[0][7] ),
	.OUT(n618));
   XOR2 U517 (.A(\mult_19_2/ab[1][5] ),
	.B(\mult_19_2/ab[0][6] ),
	.OUT(n619));
   XOR2 U518 (.A(n621),
	.B(n618),
	.OUT(n620));
   XOR2 U519 (.A(n623),
	.B(n624),
	.OUT(n622));
   XOR2 U520 (.A(\mult_19_2/ab[1][4] ),
	.B(\mult_19_2/ab[0][5] ),
	.OUT(n625));
   XOR2 U521 (.A(n627),
	.B(n619),
	.OUT(n626));
   XOR2 U522 (.A(\mult_19_2/ab[1][3] ),
	.B(\mult_19_2/ab[0][4] ),
	.OUT(n628));
   XOR2 U523 (.A(n630),
	.B(n625),
	.OUT(n629));
   XOR2 U524 (.A(n632),
	.B(n633),
	.OUT(n631));
   XOR2 U525 (.A(n635),
	.B(n636),
	.OUT(n634));
   XOR2 U526 (.A(n638),
	.B(n639),
	.OUT(n637));
   XOR2 U527 (.A(n641),
	.B(n642),
	.OUT(n640));
   XOR2 U528 (.A(n643),
	.B(n644),
	.OUT(n91));
   XOR2 U529 (.A(\mult_19_2/ab[1][2] ),
	.B(\mult_19_2/ab[0][3] ),
	.OUT(n645));
   XOR2 U530 (.A(n647),
	.B(n628),
	.OUT(n646));
   XOR2 U531 (.A(n649),
	.B(n650),
	.OUT(n648));
   XOR2 U532 (.A(n652),
	.B(n653),
	.OUT(n651));
   XOR2 U533 (.A(\mult_19_2/ab[1][1] ),
	.B(\mult_19_2/ab[0][2] ),
	.OUT(n654));
   XOR2 U534 (.A(n656),
	.B(n645),
	.OUT(n655));
   XOR2 U535 (.A(n658),
	.B(n659),
	.OUT(n657));
   XOR2 U536 (.A(n661),
	.B(n662),
	.OUT(n660));
   XOR2 U537 (.A(n664),
	.B(n665),
	.OUT(n663));
   XOR2 U538 (.A(n666),
	.B(n667),
	.OUT(n87));
   XOR2 U539 (.A(n90),
	.B(n91),
	.OUT(\mult_19_2/A1[8] ));
   XOR2 U540 (.A(n660),
	.B(n668),
	.OUT(\mult_19_2/A1[5] ));
   XOR2 U541 (.A(n657),
	.B(n669),
	.OUT(\mult_19_2/A1[3] ));
   XOR2 U542 (.A(n655),
	.B(n670),
	.OUT(\mult_19_2/A1[1] ));
   XOR2 U543 (.A(n82),
	.B(n81),
	.OUT(\mult_19_2/A1[12] ));
   XOR2 U544 (.A(n86),
	.B(n87),
	.OUT(\mult_19_2/A1[10] ));
   XOR2 U545 (.A(\mult_19/ab[1][7] ),
	.B(n672),
	.OUT(n671));
   XOR2 U546 (.A(\mult_19/ab[1][6] ),
	.B(\mult_19/ab[0][7] ),
	.OUT(n673));
   XOR2 U547 (.A(\mult_19/ab[1][5] ),
	.B(\mult_19/ab[0][6] ),
	.OUT(n674));
   XOR2 U548 (.A(n676),
	.B(n673),
	.OUT(n675));
   XOR2 U549 (.A(n678),
	.B(n679),
	.OUT(n677));
   XOR2 U550 (.A(\mult_19/ab[1][4] ),
	.B(\mult_19/ab[0][5] ),
	.OUT(n680));
   XOR2 U551 (.A(n682),
	.B(n674),
	.OUT(n681));
   XOR2 U552 (.A(\mult_19/ab[1][3] ),
	.B(\mult_19/ab[0][4] ),
	.OUT(n683));
   XOR2 U553 (.A(n685),
	.B(n680),
	.OUT(n684));
   XOR2 U554 (.A(n687),
	.B(n688),
	.OUT(n686));
   XOR2 U555 (.A(n690),
	.B(n691),
	.OUT(n689));
   XOR2 U556 (.A(n693),
	.B(n694),
	.OUT(n692));
   XOR2 U557 (.A(n696),
	.B(n697),
	.OUT(n695));
   XOR2 U558 (.A(n698),
	.B(n699),
	.OUT(n76));
   XOR2 U559 (.A(\mult_19/ab[1][2] ),
	.B(\mult_19/ab[0][3] ),
	.OUT(n700));
   XOR2 U560 (.A(n702),
	.B(n683),
	.OUT(n701));
   XOR2 U561 (.A(n704),
	.B(n705),
	.OUT(n703));
   XOR2 U562 (.A(n707),
	.B(n708),
	.OUT(n706));
   XOR2 U563 (.A(\mult_19/ab[1][1] ),
	.B(\mult_19/ab[0][2] ),
	.OUT(n709));
   XOR2 U564 (.A(n711),
	.B(n700),
	.OUT(n710));
   XOR2 U565 (.A(n713),
	.B(n714),
	.OUT(n712));
   XOR2 U566 (.A(n716),
	.B(n717),
	.OUT(n715));
   XOR2 U567 (.A(n719),
	.B(n720),
	.OUT(n718));
   XOR2 U568 (.A(n721),
	.B(n722),
	.OUT(n72));
   XOR2 U569 (.A(n75),
	.B(n76),
	.OUT(\mult_19/A1[8] ));
   XOR2 U570 (.A(n715),
	.B(n723),
	.OUT(\mult_19/A1[5] ));
   XOR2 U571 (.A(n712),
	.B(n724),
	.OUT(\mult_19/A1[3] ));
   XOR2 U572 (.A(n710),
	.B(n725),
	.OUT(\mult_19/A1[1] ));
   XOR2 U573 (.A(n67),
	.B(n66),
	.OUT(\mult_19/A1[12] ));
   XOR2 U574 (.A(n71),
	.B(n72),
	.OUT(\mult_19/A1[10] ));
   XOR2 U575 (.A(\mult_19_2/ab[1][0] ),
	.B(\mult_19_2/ab[0][1] ),
	.OUT(n726));
   XOR2 U576 (.A(\mult_19/ab[1][0] ),
	.B(\mult_19/ab[0][1] ),
	.OUT(n727));
   XOR2 U577 (.A(N17),
	.B(N1),
	.OUT(n728));
   XOR2 U578 (.A(\mult_19_3/ab[1][0] ),
	.B(\mult_19_3/ab[0][1] ),
	.OUT(n729));
   XOR2 U579 (.A(n731),
	.B(n727),
	.OUT(n730));
   XOR2 U580 (.A(\mult_21_2/ab[1][0] ),
	.B(\mult_21_2/ab[0][1] ),
	.OUT(n732));
   XOR2 U581 (.A(\mult_21/ab[1][0] ),
	.B(\mult_21/ab[0][1] ),
	.OUT(n733));
   XOR2 U582 (.A(N177),
	.B(N161),
	.OUT(n734));
   XOR2 U583 (.A(\mult_21_3/ab[1][0] ),
	.B(\mult_21_3/ab[0][1] ),
	.OUT(n735));
   XOR2 U584 (.A(n737),
	.B(n733),
	.OUT(n736));
   XOR2 U585 (.A(\mult_20_2/ab[1][0] ),
	.B(\mult_20_2/ab[0][1] ),
	.OUT(n738));
   XOR2 U586 (.A(\mult_20/ab[1][0] ),
	.B(\mult_20/ab[0][1] ),
	.OUT(n739));
   XOR2 U587 (.A(N97),
	.B(N81),
	.OUT(n740));
   XOR2 U588 (.A(\mult_20_3/ab[1][0] ),
	.B(\mult_20_3/ab[0][1] ),
	.OUT(n741));
   XOR2 U589 (.A(n743),
	.B(n739),
	.OUT(n742));
   NAND2 U590 (.A(\mult_21_3/ab[0][3] ),
	.B(\mult_21_3/ab[1][2] ),
	.OUT(n744));
   AOI21 U591 (.OUT(n745),
	.C(n747),
	.B(n746),
	.A(\mult_21_3/ab[2][2] ));
   NAND2 U592 (.A(\mult_21_3/ab[1][3] ),
	.B(\mult_21_3/ab[0][4] ),
	.OUT(n748));
   inverter U593 (.IN(\mult_21_3/ab[3][2] ),
	.OUT(n749));
   OAI21 U594 (.OUT(n750),
	.C(n751),
	.B(n749),
	.A(n745));
   NAND2 U595 (.A(\mult_21_3/ab[1][4] ),
	.B(\mult_21_3/ab[0][5] ),
	.OUT(n752));
   inverter U596 (.IN(\mult_21_3/ab[3][3] ),
	.OUT(n753));
   OAI21 U597 (.OUT(n754),
	.C(n756),
	.B(n755),
	.A(n748));
   AOI21 U598 (.OUT(n757),
	.C(n758),
	.B(\mult_21_3/ab[4][2] ),
	.A(n750));
   NAND2 U599 (.A(\mult_21_3/ab[1][5] ),
	.B(\mult_21_3/ab[0][6] ),
	.OUT(n759));
   inverter U600 (.IN(\mult_21_3/ab[3][4] ),
	.OUT(n760));
   OAI21 U601 (.OUT(n761),
	.C(n763),
	.B(n762),
	.A(n752));
   AOI21 U602 (.OUT(n764),
	.C(n765),
	.B(\mult_21_3/ab[3][3] ),
	.A(n754));
   inverter U603 (.IN(\mult_21_3/ab[5][2] ),
	.OUT(n766));
   OAI21 U604 (.OUT(n767),
	.C(n768),
	.B(n766),
	.A(n757));
   NAND2 U605 (.A(\mult_21_3/ab[1][6] ),
	.B(\mult_21_3/ab[0][7] ),
	.OUT(n769));
   OAI21 U606 (.OUT(n770),
	.C(n772),
	.B(n771),
	.A(n759));
   inverter U607 (.IN(\mult_21_3/ab[4][4] ),
	.OUT(n773));
   AOI21 U608 (.OUT(n774),
	.C(n775),
	.B(\mult_21_3/ab[3][4] ),
	.A(n761));
   OAI21 U609 (.OUT(n776),
	.C(n778),
	.B(n777),
	.A(n764));
   AOI21 U610 (.OUT(n779),
	.C(n780),
	.B(\mult_21_3/ab[6][2] ),
	.A(n767));
   inverter U611 (.IN(\mult_21_3/ab[3][6] ),
	.OUT(n781));
   inverter U612 (.IN(\mult_21_3/ab[2][7] ),
	.OUT(n782));
   OAI21 U613 (.OUT(n783),
	.C(n786),
	.B(n785),
	.A(n784));
   inverter U614 (.IN(\mult_21_3/ab[5][4] ),
	.OUT(n787));
   AOI21 U615 (.OUT(n788),
	.C(n790),
	.B(\mult_21_3/ab[4][4] ),
	.A(n789));
   AOI21 U616 (.OUT(n791),
	.C(n792),
	.B(\mult_21_3/ab[5][3] ),
	.A(n776));
   inverter U617 (.IN(\mult_21_3/ab[4][6] ),
	.OUT(n793));
   inverter U618 (.IN(\mult_21_3/ab[3][7] ),
	.OUT(n794));
   AOI21 U619 (.OUT(n795),
	.C(n796),
	.B(\mult_21_3/ab[4][5] ),
	.A(n783));
   OAI21 U620 (.OUT(n797),
	.C(n798),
	.B(n787),
	.A(n788));
   OAI21 U621 (.OUT(n799),
	.C(n801),
	.B(n800),
	.A(n791));
   NAND2 U622 (.A(\mult_21_3/ab[0][2] ),
	.B(\mult_21_3/ab[1][1] ),
	.OUT(n802));
   OAI21 U623 (.OUT(n803),
	.C(n805),
	.B(n802),
	.A(n804));
   inverter U624 (.IN(\mult_21_3/ab[3][1] ),
	.OUT(n806));
   AOI21 U625 (.OUT(n807),
	.C(n808),
	.B(\mult_21_3/ab[3][1] ),
	.A(n803));
   OAI21 U626 (.OUT(n809),
	.C(n811),
	.B(n810),
	.A(n807));
   AOI21 U627 (.OUT(n812),
	.C(n813),
	.B(\mult_21_3/ab[5][1] ),
	.A(n809));
   inverter U628 (.IN(\mult_21_3/ab[6][1] ),
	.OUT(n814));
   OAI21 U629 (.OUT(n815),
	.C(n816),
	.B(n814),
	.A(n812));
   NAND2 U630 (.A(\mult_21_3/ab[0][1] ),
	.B(\mult_21_3/ab[1][0] ),
	.OUT(n817));
   AOI21 U631 (.OUT(n818),
	.C(n820),
	.B(n819),
	.A(\mult_21_3/ab[2][0] ));
   inverter U632 (.IN(\mult_21_3/ab[3][0] ),
	.OUT(n821));
   OAI21 U633 (.OUT(n822),
	.C(n823),
	.B(n821),
	.A(n818));
   AOI21 U634 (.OUT(n824),
	.C(n825),
	.B(\mult_21_3/ab[4][0] ),
	.A(n822));
   inverter U635 (.IN(\mult_21_3/ab[5][0] ),
	.OUT(n826));
   OAI21 U636 (.OUT(n827),
	.C(n828),
	.B(n826),
	.A(n824));
   AOI21 U637 (.OUT(n829),
	.C(n830),
	.B(\mult_21_3/ab[6][0] ),
	.A(n827));
   inverter U638 (.IN(\mult_21_3/ab[7][0] ),
	.OUT(n831));
   inverter U639 (.IN(\mult_21_3/ab[4][7] ),
	.OUT(n832));
   inverter U640 (.IN(\mult_21_3/ab[5][6] ),
	.OUT(n833));
   inverter U641 (.IN(\mult_21_3/ab[5][7] ),
	.OUT(n834));
   inverter U642 (.IN(\mult_21_3/ab[6][6] ),
	.OUT(n835));
   inverter U643 (.IN(\mult_21_3/ab[7][7] ),
	.OUT(n187));
   AOI21 U644 (.OUT(n836),
	.C(n838),
	.B(\mult_21_3/ab[5][5] ),
	.A(n837));
   inverter U645 (.IN(\mult_21_3/ab[6][5] ),
	.OUT(n839));
   OAI21 U646 (.OUT(n840),
	.C(n841),
	.B(n839),
	.A(n836));
   AOI21 U647 (.OUT(n842),
	.C(n843),
	.B(\mult_21_3/ab[6][4] ),
	.A(n797));
   NAND2 U648 (.A(\mult_21_2/ab[0][3] ),
	.B(\mult_21_2/ab[1][2] ),
	.OUT(n844));
   AOI21 U649 (.OUT(n845),
	.C(n847),
	.B(n846),
	.A(\mult_21_2/ab[2][2] ));
   NAND2 U650 (.A(\mult_21_2/ab[1][3] ),
	.B(\mult_21_2/ab[0][4] ),
	.OUT(n848));
   inverter U651 (.IN(\mult_21_2/ab[3][2] ),
	.OUT(n849));
   OAI21 U652 (.OUT(n850),
	.C(n851),
	.B(n849),
	.A(n845));
   NAND2 U653 (.A(\mult_21_2/ab[1][4] ),
	.B(\mult_21_2/ab[0][5] ),
	.OUT(n852));
   inverter U654 (.IN(\mult_21_2/ab[3][3] ),
	.OUT(n853));
   OAI21 U655 (.OUT(n854),
	.C(n856),
	.B(n855),
	.A(n848));
   AOI21 U656 (.OUT(n857),
	.C(n858),
	.B(\mult_21_2/ab[4][2] ),
	.A(n850));
   NAND2 U657 (.A(\mult_21_2/ab[1][5] ),
	.B(\mult_21_2/ab[0][6] ),
	.OUT(n859));
   inverter U658 (.IN(\mult_21_2/ab[3][4] ),
	.OUT(n860));
   OAI21 U659 (.OUT(n861),
	.C(n863),
	.B(n862),
	.A(n852));
   AOI21 U660 (.OUT(n864),
	.C(n865),
	.B(\mult_21_2/ab[3][3] ),
	.A(n854));
   inverter U661 (.IN(\mult_21_2/ab[5][2] ),
	.OUT(n866));
   OAI21 U662 (.OUT(n867),
	.C(n868),
	.B(n866),
	.A(n857));
   NAND2 U663 (.A(\mult_21_2/ab[1][6] ),
	.B(\mult_21_2/ab[0][7] ),
	.OUT(n869));
   OAI21 U664 (.OUT(n870),
	.C(n872),
	.B(n871),
	.A(n859));
   inverter U665 (.IN(\mult_21_2/ab[4][4] ),
	.OUT(n873));
   AOI21 U666 (.OUT(n874),
	.C(n875),
	.B(\mult_21_2/ab[3][4] ),
	.A(n861));
   OAI21 U667 (.OUT(n876),
	.C(n878),
	.B(n877),
	.A(n864));
   AOI21 U668 (.OUT(n879),
	.C(n880),
	.B(\mult_21_2/ab[6][2] ),
	.A(n867));
   inverter U669 (.IN(\mult_21_2/ab[3][6] ),
	.OUT(n881));
   inverter U670 (.IN(\mult_21_2/ab[2][7] ),
	.OUT(n882));
   OAI21 U671 (.OUT(n883),
	.C(n886),
	.B(n885),
	.A(n884));
   inverter U672 (.IN(\mult_21_2/ab[5][4] ),
	.OUT(n887));
   AOI21 U673 (.OUT(n888),
	.C(n890),
	.B(\mult_21_2/ab[4][4] ),
	.A(n889));
   AOI21 U674 (.OUT(n891),
	.C(n892),
	.B(\mult_21_2/ab[5][3] ),
	.A(n876));
   inverter U675 (.IN(\mult_21_2/ab[4][6] ),
	.OUT(n893));
   inverter U676 (.IN(\mult_21_2/ab[3][7] ),
	.OUT(n894));
   AOI21 U677 (.OUT(n895),
	.C(n896),
	.B(\mult_21_2/ab[4][5] ),
	.A(n883));
   OAI21 U678 (.OUT(n897),
	.C(n898),
	.B(n887),
	.A(n888));
   OAI21 U679 (.OUT(n899),
	.C(n901),
	.B(n900),
	.A(n891));
   NAND2 U680 (.A(\mult_21_2/ab[0][2] ),
	.B(\mult_21_2/ab[1][1] ),
	.OUT(n902));
   OAI21 U681 (.OUT(n903),
	.C(n905),
	.B(n902),
	.A(n904));
   inverter U682 (.IN(\mult_21_2/ab[3][1] ),
	.OUT(n906));
   AOI21 U683 (.OUT(n907),
	.C(n908),
	.B(\mult_21_2/ab[3][1] ),
	.A(n903));
   OAI21 U684 (.OUT(n909),
	.C(n911),
	.B(n910),
	.A(n907));
   AOI21 U685 (.OUT(n912),
	.C(n913),
	.B(\mult_21_2/ab[5][1] ),
	.A(n909));
   inverter U686 (.IN(\mult_21_2/ab[6][1] ),
	.OUT(n914));
   OAI21 U687 (.OUT(n915),
	.C(n916),
	.B(n914),
	.A(n912));
   NAND2 U688 (.A(\mult_21_2/ab[0][1] ),
	.B(\mult_21_2/ab[1][0] ),
	.OUT(n917));
   AOI21 U689 (.OUT(n918),
	.C(n920),
	.B(n919),
	.A(\mult_21_2/ab[2][0] ));
   inverter U690 (.IN(\mult_21_2/ab[3][0] ),
	.OUT(n921));
   OAI21 U691 (.OUT(n922),
	.C(n923),
	.B(n921),
	.A(n918));
   AOI21 U692 (.OUT(n924),
	.C(n925),
	.B(\mult_21_2/ab[4][0] ),
	.A(n922));
   inverter U693 (.IN(\mult_21_2/ab[5][0] ),
	.OUT(n926));
   OAI21 U694 (.OUT(n927),
	.C(n928),
	.B(n926),
	.A(n924));
   AOI21 U695 (.OUT(n929),
	.C(n930),
	.B(\mult_21_2/ab[6][0] ),
	.A(n927));
   inverter U696 (.IN(\mult_21_2/ab[7][0] ),
	.OUT(n931));
   inverter U697 (.IN(\mult_21_2/ab[4][7] ),
	.OUT(n932));
   inverter U698 (.IN(\mult_21_2/ab[5][6] ),
	.OUT(n933));
   inverter U699 (.IN(\mult_21_2/ab[5][7] ),
	.OUT(n934));
   inverter U700 (.IN(\mult_21_2/ab[6][6] ),
	.OUT(n935));
   inverter U701 (.IN(\mult_21_2/ab[7][7] ),
	.OUT(n172));
   AOI21 U702 (.OUT(n936),
	.C(n938),
	.B(\mult_21_2/ab[5][5] ),
	.A(n937));
   inverter U703 (.IN(\mult_21_2/ab[6][5] ),
	.OUT(n939));
   OAI21 U704 (.OUT(n940),
	.C(n941),
	.B(n939),
	.A(n936));
   AOI21 U705 (.OUT(n942),
	.C(n943),
	.B(\mult_21_2/ab[6][4] ),
	.A(n897));
   NAND2 U706 (.A(\mult_21/ab[0][3] ),
	.B(\mult_21/ab[1][2] ),
	.OUT(n944));
   AOI21 U707 (.OUT(n945),
	.C(n947),
	.B(n946),
	.A(\mult_21/ab[2][2] ));
   NAND2 U708 (.A(\mult_21/ab[1][3] ),
	.B(\mult_21/ab[0][4] ),
	.OUT(n948));
   inverter U709 (.IN(\mult_21/ab[3][2] ),
	.OUT(n949));
   OAI21 U710 (.OUT(n950),
	.C(n951),
	.B(n949),
	.A(n945));
   NAND2 U711 (.A(\mult_21/ab[1][4] ),
	.B(\mult_21/ab[0][5] ),
	.OUT(n952));
   inverter U712 (.IN(\mult_21/ab[3][3] ),
	.OUT(n953));
   OAI21 U713 (.OUT(n954),
	.C(n956),
	.B(n955),
	.A(n948));
   AOI21 U714 (.OUT(n957),
	.C(n958),
	.B(\mult_21/ab[4][2] ),
	.A(n950));
   NAND2 U715 (.A(\mult_21/ab[1][5] ),
	.B(\mult_21/ab[0][6] ),
	.OUT(n959));
   inverter U716 (.IN(\mult_21/ab[3][4] ),
	.OUT(n960));
   OAI21 U717 (.OUT(n961),
	.C(n963),
	.B(n962),
	.A(n952));
   AOI21 U718 (.OUT(n964),
	.C(n965),
	.B(\mult_21/ab[3][3] ),
	.A(n954));
   inverter U719 (.IN(\mult_21/ab[5][2] ),
	.OUT(n966));
   OAI21 U720 (.OUT(n967),
	.C(n968),
	.B(n966),
	.A(n957));
   NAND2 U721 (.A(\mult_21/ab[1][6] ),
	.B(\mult_21/ab[0][7] ),
	.OUT(n969));
   OAI21 U722 (.OUT(n970),
	.C(n972),
	.B(n971),
	.A(n959));
   inverter U723 (.IN(\mult_21/ab[4][4] ),
	.OUT(n973));
   AOI21 U724 (.OUT(n974),
	.C(n975),
	.B(\mult_21/ab[3][4] ),
	.A(n961));
   OAI21 U725 (.OUT(n976),
	.C(n978),
	.B(n977),
	.A(n964));
   AOI21 U726 (.OUT(n979),
	.C(n980),
	.B(\mult_21/ab[6][2] ),
	.A(n967));
   inverter U727 (.IN(\mult_21/ab[3][6] ),
	.OUT(n981));
   inverter U728 (.IN(\mult_21/ab[2][7] ),
	.OUT(n982));
   OAI21 U729 (.OUT(n983),
	.C(n986),
	.B(n985),
	.A(n984));
   inverter U730 (.IN(\mult_21/ab[5][4] ),
	.OUT(n987));
   AOI21 U731 (.OUT(n988),
	.C(n990),
	.B(\mult_21/ab[4][4] ),
	.A(n989));
   AOI21 U732 (.OUT(n991),
	.C(n992),
	.B(\mult_21/ab[5][3] ),
	.A(n976));
   inverter U733 (.IN(\mult_21/ab[4][6] ),
	.OUT(n993));
   inverter U734 (.IN(\mult_21/ab[3][7] ),
	.OUT(n994));
   AOI21 U735 (.OUT(n995),
	.C(n996),
	.B(\mult_21/ab[4][5] ),
	.A(n983));
   OAI21 U736 (.OUT(n997),
	.C(n998),
	.B(n987),
	.A(n988));
   OAI21 U737 (.OUT(n999),
	.C(n1001),
	.B(n1000),
	.A(n991));
   NAND2 U738 (.A(\mult_21/ab[0][2] ),
	.B(\mult_21/ab[1][1] ),
	.OUT(n1002));
   OAI21 U739 (.OUT(n1003),
	.C(n1005),
	.B(n1002),
	.A(n1004));
   inverter U740 (.IN(\mult_21/ab[3][1] ),
	.OUT(n1006));
   AOI21 U741 (.OUT(n1007),
	.C(n1008),
	.B(\mult_21/ab[3][1] ),
	.A(n1003));
   OAI21 U742 (.OUT(n1009),
	.C(n1011),
	.B(n1010),
	.A(n1007));
   AOI21 U743 (.OUT(n1012),
	.C(n1013),
	.B(\mult_21/ab[5][1] ),
	.A(n1009));
   inverter U744 (.IN(\mult_21/ab[6][1] ),
	.OUT(n1014));
   OAI21 U745 (.OUT(n1015),
	.C(n1016),
	.B(n1014),
	.A(n1012));
   NAND2 U746 (.A(\mult_21/ab[0][1] ),
	.B(\mult_21/ab[1][0] ),
	.OUT(n1017));
   AOI21 U747 (.OUT(n1018),
	.C(n1020),
	.B(n1019),
	.A(\mult_21/ab[2][0] ));
   inverter U748 (.IN(\mult_21/ab[3][0] ),
	.OUT(n1021));
   OAI21 U749 (.OUT(n1022),
	.C(n1023),
	.B(n1021),
	.A(n1018));
   AOI21 U750 (.OUT(n1024),
	.C(n1025),
	.B(\mult_21/ab[4][0] ),
	.A(n1022));
   inverter U751 (.IN(\mult_21/ab[5][0] ),
	.OUT(n1026));
   OAI21 U752 (.OUT(n1027),
	.C(n1028),
	.B(n1026),
	.A(n1024));
   AOI21 U753 (.OUT(n1029),
	.C(n1030),
	.B(\mult_21/ab[6][0] ),
	.A(n1027));
   inverter U754 (.IN(\mult_21/ab[7][0] ),
	.OUT(n1031));
   inverter U755 (.IN(\mult_21/ab[4][7] ),
	.OUT(n1032));
   inverter U756 (.IN(\mult_21/ab[5][6] ),
	.OUT(n1033));
   inverter U757 (.IN(\mult_21/ab[5][7] ),
	.OUT(n1034));
   inverter U758 (.IN(\mult_21/ab[6][6] ),
	.OUT(n1035));
   inverter U759 (.IN(\mult_21/ab[7][7] ),
	.OUT(n157));
   AOI21 U760 (.OUT(n1036),
	.C(n1038),
	.B(\mult_21/ab[5][5] ),
	.A(n1037));
   inverter U761 (.IN(\mult_21/ab[6][5] ),
	.OUT(n1039));
   OAI21 U762 (.OUT(n1040),
	.C(n1041),
	.B(n1039),
	.A(n1036));
   AOI21 U763 (.OUT(n1042),
	.C(n1043),
	.B(\mult_21/ab[6][4] ),
	.A(n997));
   NAND2 U764 (.A(\mult_20_3/ab[0][3] ),
	.B(\mult_20_3/ab[1][2] ),
	.OUT(n1044));
   AOI21 U765 (.OUT(n1045),
	.C(n1047),
	.B(n1046),
	.A(\mult_20_3/ab[2][2] ));
   NAND2 U766 (.A(\mult_20_3/ab[1][3] ),
	.B(\mult_20_3/ab[0][4] ),
	.OUT(n1048));
   inverter U767 (.IN(\mult_20_3/ab[3][2] ),
	.OUT(n1049));
   OAI21 U768 (.OUT(n1050),
	.C(n1051),
	.B(n1049),
	.A(n1045));
   NAND2 U769 (.A(\mult_20_3/ab[1][4] ),
	.B(\mult_20_3/ab[0][5] ),
	.OUT(n1052));
   inverter U770 (.IN(\mult_20_3/ab[3][3] ),
	.OUT(n1053));
   OAI21 U771 (.OUT(n1054),
	.C(n1056),
	.B(n1055),
	.A(n1048));
   AOI21 U772 (.OUT(n1057),
	.C(n1058),
	.B(\mult_20_3/ab[4][2] ),
	.A(n1050));
   NAND2 U773 (.A(\mult_20_3/ab[1][5] ),
	.B(\mult_20_3/ab[0][6] ),
	.OUT(n1059));
   inverter U774 (.IN(\mult_20_3/ab[3][4] ),
	.OUT(n1060));
   OAI21 U775 (.OUT(n1061),
	.C(n1063),
	.B(n1062),
	.A(n1052));
   AOI21 U776 (.OUT(n1064),
	.C(n1065),
	.B(\mult_20_3/ab[3][3] ),
	.A(n1054));
   inverter U777 (.IN(\mult_20_3/ab[5][2] ),
	.OUT(n1066));
   OAI21 U778 (.OUT(n1067),
	.C(n1068),
	.B(n1066),
	.A(n1057));
   NAND2 U779 (.A(\mult_20_3/ab[1][6] ),
	.B(\mult_20_3/ab[0][7] ),
	.OUT(n1069));
   OAI21 U780 (.OUT(n1070),
	.C(n1072),
	.B(n1071),
	.A(n1059));
   inverter U781 (.IN(\mult_20_3/ab[4][4] ),
	.OUT(n1073));
   AOI21 U782 (.OUT(n1074),
	.C(n1075),
	.B(\mult_20_3/ab[3][4] ),
	.A(n1061));
   OAI21 U783 (.OUT(n1076),
	.C(n1078),
	.B(n1077),
	.A(n1064));
   AOI21 U784 (.OUT(n1079),
	.C(n1080),
	.B(\mult_20_3/ab[6][2] ),
	.A(n1067));
   inverter U785 (.IN(\mult_20_3/ab[3][6] ),
	.OUT(n1081));
   inverter U786 (.IN(\mult_20_3/ab[2][7] ),
	.OUT(n1082));
   OAI21 U787 (.OUT(n1083),
	.C(n1086),
	.B(n1085),
	.A(n1084));
   inverter U788 (.IN(\mult_20_3/ab[5][4] ),
	.OUT(n1087));
   AOI21 U789 (.OUT(n1088),
	.C(n1090),
	.B(\mult_20_3/ab[4][4] ),
	.A(n1089));
   AOI21 U790 (.OUT(n1091),
	.C(n1092),
	.B(\mult_20_3/ab[5][3] ),
	.A(n1076));
   inverter U791 (.IN(\mult_20_3/ab[4][6] ),
	.OUT(n1093));
   inverter U792 (.IN(\mult_20_3/ab[3][7] ),
	.OUT(n1094));
   AOI21 U793 (.OUT(n1095),
	.C(n1096),
	.B(\mult_20_3/ab[4][5] ),
	.A(n1083));
   OAI21 U794 (.OUT(n1097),
	.C(n1098),
	.B(n1087),
	.A(n1088));
   OAI21 U795 (.OUT(n1099),
	.C(n1101),
	.B(n1100),
	.A(n1091));
   NAND2 U796 (.A(\mult_20_3/ab[0][2] ),
	.B(\mult_20_3/ab[1][1] ),
	.OUT(n1102));
   OAI21 U797 (.OUT(n1103),
	.C(n1105),
	.B(n1102),
	.A(n1104));
   inverter U798 (.IN(\mult_20_3/ab[3][1] ),
	.OUT(n1106));
   AOI21 U799 (.OUT(n1107),
	.C(n1108),
	.B(\mult_20_3/ab[3][1] ),
	.A(n1103));
   OAI21 U800 (.OUT(n1109),
	.C(n1111),
	.B(n1110),
	.A(n1107));
   AOI21 U801 (.OUT(n1112),
	.C(n1113),
	.B(\mult_20_3/ab[5][1] ),
	.A(n1109));
   inverter U802 (.IN(\mult_20_3/ab[6][1] ),
	.OUT(n1114));
   OAI21 U803 (.OUT(n1115),
	.C(n1116),
	.B(n1114),
	.A(n1112));
   NAND2 U804 (.A(\mult_20_3/ab[0][1] ),
	.B(\mult_20_3/ab[1][0] ),
	.OUT(n1117));
   AOI21 U805 (.OUT(n1118),
	.C(n1120),
	.B(n1119),
	.A(\mult_20_3/ab[2][0] ));
   inverter U806 (.IN(\mult_20_3/ab[3][0] ),
	.OUT(n1121));
   OAI21 U807 (.OUT(n1122),
	.C(n1123),
	.B(n1121),
	.A(n1118));
   AOI21 U808 (.OUT(n1124),
	.C(n1125),
	.B(\mult_20_3/ab[4][0] ),
	.A(n1122));
   inverter U809 (.IN(\mult_20_3/ab[5][0] ),
	.OUT(n1126));
   OAI21 U810 (.OUT(n1127),
	.C(n1128),
	.B(n1126),
	.A(n1124));
   AOI21 U811 (.OUT(n1129),
	.C(n1130),
	.B(\mult_20_3/ab[6][0] ),
	.A(n1127));
   inverter U812 (.IN(\mult_20_3/ab[7][0] ),
	.OUT(n1131));
   inverter U813 (.IN(\mult_20_3/ab[4][7] ),
	.OUT(n1132));
   inverter U814 (.IN(\mult_20_3/ab[5][6] ),
	.OUT(n1133));
   inverter U815 (.IN(\mult_20_3/ab[5][7] ),
	.OUT(n1134));
   inverter U816 (.IN(\mult_20_3/ab[6][6] ),
	.OUT(n1135));
   inverter U817 (.IN(\mult_20_3/ab[7][7] ),
	.OUT(n142));
   AOI21 U818 (.OUT(n1136),
	.C(n1138),
	.B(\mult_20_3/ab[5][5] ),
	.A(n1137));
   inverter U819 (.IN(\mult_20_3/ab[6][5] ),
	.OUT(n1139));
   OAI21 U820 (.OUT(n1140),
	.C(n1141),
	.B(n1139),
	.A(n1136));
   AOI21 U821 (.OUT(n1142),
	.C(n1143),
	.B(\mult_20_3/ab[6][4] ),
	.A(n1097));
   NAND2 U822 (.A(\mult_20_2/ab[0][3] ),
	.B(\mult_20_2/ab[1][2] ),
	.OUT(n1144));
   AOI21 U823 (.OUT(n1145),
	.C(n1147),
	.B(n1146),
	.A(\mult_20_2/ab[2][2] ));
   NAND2 U824 (.A(\mult_20_2/ab[1][3] ),
	.B(\mult_20_2/ab[0][4] ),
	.OUT(n1148));
   inverter U825 (.IN(\mult_20_2/ab[3][2] ),
	.OUT(n1149));
   OAI21 U826 (.OUT(n1150),
	.C(n1151),
	.B(n1149),
	.A(n1145));
   NAND2 U827 (.A(\mult_20_2/ab[1][4] ),
	.B(\mult_20_2/ab[0][5] ),
	.OUT(n1152));
   inverter U828 (.IN(\mult_20_2/ab[3][3] ),
	.OUT(n1153));
   OAI21 U829 (.OUT(n1154),
	.C(n1156),
	.B(n1155),
	.A(n1148));
   AOI21 U830 (.OUT(n1157),
	.C(n1158),
	.B(\mult_20_2/ab[4][2] ),
	.A(n1150));
   NAND2 U831 (.A(\mult_20_2/ab[1][5] ),
	.B(\mult_20_2/ab[0][6] ),
	.OUT(n1159));
   inverter U832 (.IN(\mult_20_2/ab[3][4] ),
	.OUT(n1160));
   OAI21 U833 (.OUT(n1161),
	.C(n1163),
	.B(n1162),
	.A(n1152));
   AOI21 U834 (.OUT(n1164),
	.C(n1165),
	.B(\mult_20_2/ab[3][3] ),
	.A(n1154));
   inverter U835 (.IN(\mult_20_2/ab[5][2] ),
	.OUT(n1166));
   OAI21 U836 (.OUT(n1167),
	.C(n1168),
	.B(n1166),
	.A(n1157));
   NAND2 U837 (.A(\mult_20_2/ab[1][6] ),
	.B(\mult_20_2/ab[0][7] ),
	.OUT(n1169));
   OAI21 U838 (.OUT(n1170),
	.C(n1172),
	.B(n1171),
	.A(n1159));
   inverter U839 (.IN(\mult_20_2/ab[4][4] ),
	.OUT(n1173));
   AOI21 U840 (.OUT(n1174),
	.C(n1175),
	.B(\mult_20_2/ab[3][4] ),
	.A(n1161));
   OAI21 U841 (.OUT(n1176),
	.C(n1178),
	.B(n1177),
	.A(n1164));
   AOI21 U842 (.OUT(n1179),
	.C(n1180),
	.B(\mult_20_2/ab[6][2] ),
	.A(n1167));
   inverter U843 (.IN(\mult_20_2/ab[3][6] ),
	.OUT(n1181));
   inverter U844 (.IN(\mult_20_2/ab[2][7] ),
	.OUT(n1182));
   OAI21 U845 (.OUT(n1183),
	.C(n1186),
	.B(n1185),
	.A(n1184));
   inverter U846 (.IN(\mult_20_2/ab[5][4] ),
	.OUT(n1187));
   AOI21 U847 (.OUT(n1188),
	.C(n1190),
	.B(\mult_20_2/ab[4][4] ),
	.A(n1189));
   AOI21 U848 (.OUT(n1191),
	.C(n1192),
	.B(\mult_20_2/ab[5][3] ),
	.A(n1176));
   inverter U849 (.IN(\mult_20_2/ab[4][6] ),
	.OUT(n1193));
   inverter U850 (.IN(\mult_20_2/ab[3][7] ),
	.OUT(n1194));
   AOI21 U851 (.OUT(n1195),
	.C(n1196),
	.B(\mult_20_2/ab[4][5] ),
	.A(n1183));
   OAI21 U852 (.OUT(n1197),
	.C(n1198),
	.B(n1187),
	.A(n1188));
   OAI21 U853 (.OUT(n1199),
	.C(n1201),
	.B(n1200),
	.A(n1191));
   NAND2 U854 (.A(\mult_20_2/ab[0][2] ),
	.B(\mult_20_2/ab[1][1] ),
	.OUT(n1202));
   OAI21 U855 (.OUT(n1203),
	.C(n1205),
	.B(n1202),
	.A(n1204));
   inverter U856 (.IN(\mult_20_2/ab[3][1] ),
	.OUT(n1206));
   AOI21 U857 (.OUT(n1207),
	.C(n1208),
	.B(\mult_20_2/ab[3][1] ),
	.A(n1203));
   OAI21 U858 (.OUT(n1209),
	.C(n1211),
	.B(n1210),
	.A(n1207));
   AOI21 U859 (.OUT(n1212),
	.C(n1213),
	.B(\mult_20_2/ab[5][1] ),
	.A(n1209));
   inverter U860 (.IN(\mult_20_2/ab[6][1] ),
	.OUT(n1214));
   OAI21 U861 (.OUT(n1215),
	.C(n1216),
	.B(n1214),
	.A(n1212));
   NAND2 U862 (.A(\mult_20_2/ab[0][1] ),
	.B(\mult_20_2/ab[1][0] ),
	.OUT(n1217));
   AOI21 U863 (.OUT(n1218),
	.C(n1220),
	.B(n1219),
	.A(\mult_20_2/ab[2][0] ));
   inverter U864 (.IN(\mult_20_2/ab[3][0] ),
	.OUT(n1221));
   OAI21 U865 (.OUT(n1222),
	.C(n1223),
	.B(n1221),
	.A(n1218));
   AOI21 U866 (.OUT(n1224),
	.C(n1225),
	.B(\mult_20_2/ab[4][0] ),
	.A(n1222));
   inverter U867 (.IN(\mult_20_2/ab[5][0] ),
	.OUT(n1226));
   OAI21 U868 (.OUT(n1227),
	.C(n1228),
	.B(n1226),
	.A(n1224));
   AOI21 U869 (.OUT(n1229),
	.C(n1230),
	.B(\mult_20_2/ab[6][0] ),
	.A(n1227));
   inverter U870 (.IN(\mult_20_2/ab[7][0] ),
	.OUT(n1231));
   inverter U871 (.IN(\mult_20_2/ab[4][7] ),
	.OUT(n1232));
   inverter U872 (.IN(\mult_20_2/ab[5][6] ),
	.OUT(n1233));
   inverter U873 (.IN(\mult_20_2/ab[5][7] ),
	.OUT(n1234));
   inverter U874 (.IN(\mult_20_2/ab[6][6] ),
	.OUT(n1235));
   inverter U875 (.IN(\mult_20_2/ab[7][7] ),
	.OUT(n127));
   AOI21 U876 (.OUT(n1236),
	.C(n1238),
	.B(\mult_20_2/ab[5][5] ),
	.A(n1237));
   inverter U877 (.IN(\mult_20_2/ab[6][5] ),
	.OUT(n1239));
   OAI21 U878 (.OUT(n1240),
	.C(n1241),
	.B(n1239),
	.A(n1236));
   AOI21 U879 (.OUT(n1242),
	.C(n1243),
	.B(\mult_20_2/ab[6][4] ),
	.A(n1197));
   NAND2 U880 (.A(\mult_20/ab[0][3] ),
	.B(\mult_20/ab[1][2] ),
	.OUT(n1244));
   AOI21 U881 (.OUT(n1245),
	.C(n1247),
	.B(n1246),
	.A(\mult_20/ab[2][2] ));
   NAND2 U882 (.A(\mult_20/ab[1][3] ),
	.B(\mult_20/ab[0][4] ),
	.OUT(n1248));
   inverter U883 (.IN(\mult_20/ab[3][2] ),
	.OUT(n1249));
   OAI21 U884 (.OUT(n1250),
	.C(n1251),
	.B(n1249),
	.A(n1245));
   NAND2 U885 (.A(\mult_20/ab[1][4] ),
	.B(\mult_20/ab[0][5] ),
	.OUT(n1252));
   inverter U886 (.IN(\mult_20/ab[3][3] ),
	.OUT(n1253));
   OAI21 U887 (.OUT(n1254),
	.C(n1256),
	.B(n1255),
	.A(n1248));
   AOI21 U888 (.OUT(n1257),
	.C(n1258),
	.B(\mult_20/ab[4][2] ),
	.A(n1250));
   NAND2 U889 (.A(\mult_20/ab[1][5] ),
	.B(\mult_20/ab[0][6] ),
	.OUT(n1259));
   inverter U890 (.IN(\mult_20/ab[3][4] ),
	.OUT(n1260));
   OAI21 U891 (.OUT(n1261),
	.C(n1263),
	.B(n1262),
	.A(n1252));
   AOI21 U892 (.OUT(n1264),
	.C(n1265),
	.B(\mult_20/ab[3][3] ),
	.A(n1254));
   inverter U893 (.IN(\mult_20/ab[5][2] ),
	.OUT(n1266));
   OAI21 U894 (.OUT(n1267),
	.C(n1268),
	.B(n1266),
	.A(n1257));
   NAND2 U895 (.A(\mult_20/ab[1][6] ),
	.B(\mult_20/ab[0][7] ),
	.OUT(n1269));
   OAI21 U896 (.OUT(n1270),
	.C(n1272),
	.B(n1271),
	.A(n1259));
   inverter U897 (.IN(\mult_20/ab[4][4] ),
	.OUT(n1273));
   AOI21 U898 (.OUT(n1274),
	.C(n1275),
	.B(\mult_20/ab[3][4] ),
	.A(n1261));
   OAI21 U899 (.OUT(n1276),
	.C(n1278),
	.B(n1277),
	.A(n1264));
   AOI21 U900 (.OUT(n1279),
	.C(n1280),
	.B(\mult_20/ab[6][2] ),
	.A(n1267));
   inverter U901 (.IN(\mult_20/ab[3][6] ),
	.OUT(n1281));
   inverter U902 (.IN(\mult_20/ab[2][7] ),
	.OUT(n1282));
   OAI21 U903 (.OUT(n1283),
	.C(n1286),
	.B(n1285),
	.A(n1284));
   inverter U904 (.IN(\mult_20/ab[5][4] ),
	.OUT(n1287));
   AOI21 U905 (.OUT(n1288),
	.C(n1290),
	.B(\mult_20/ab[4][4] ),
	.A(n1289));
   AOI21 U906 (.OUT(n1291),
	.C(n1292),
	.B(\mult_20/ab[5][3] ),
	.A(n1276));
   inverter U907 (.IN(\mult_20/ab[4][6] ),
	.OUT(n1293));
   inverter U908 (.IN(\mult_20/ab[3][7] ),
	.OUT(n1294));
   AOI21 U909 (.OUT(n1295),
	.C(n1296),
	.B(\mult_20/ab[4][5] ),
	.A(n1283));
   OAI21 U910 (.OUT(n1297),
	.C(n1298),
	.B(n1287),
	.A(n1288));
   OAI21 U911 (.OUT(n1299),
	.C(n1301),
	.B(n1300),
	.A(n1291));
   NAND2 U912 (.A(\mult_20/ab[0][2] ),
	.B(\mult_20/ab[1][1] ),
	.OUT(n1302));
   OAI21 U913 (.OUT(n1303),
	.C(n1305),
	.B(n1302),
	.A(n1304));
   inverter U914 (.IN(\mult_20/ab[3][1] ),
	.OUT(n1306));
   AOI21 U915 (.OUT(n1307),
	.C(n1308),
	.B(\mult_20/ab[3][1] ),
	.A(n1303));
   OAI21 U916 (.OUT(n1309),
	.C(n1311),
	.B(n1310),
	.A(n1307));
   AOI21 U917 (.OUT(n1312),
	.C(n1313),
	.B(\mult_20/ab[5][1] ),
	.A(n1309));
   inverter U918 (.IN(\mult_20/ab[6][1] ),
	.OUT(n1314));
   OAI21 U919 (.OUT(n1315),
	.C(n1316),
	.B(n1314),
	.A(n1312));
   NAND2 U920 (.A(\mult_20/ab[0][1] ),
	.B(\mult_20/ab[1][0] ),
	.OUT(n1317));
   AOI21 U921 (.OUT(n1318),
	.C(n1320),
	.B(n1319),
	.A(\mult_20/ab[2][0] ));
   inverter U922 (.IN(\mult_20/ab[3][0] ),
	.OUT(n1321));
   OAI21 U923 (.OUT(n1322),
	.C(n1323),
	.B(n1321),
	.A(n1318));
   AOI21 U924 (.OUT(n1324),
	.C(n1325),
	.B(\mult_20/ab[4][0] ),
	.A(n1322));
   inverter U925 (.IN(\mult_20/ab[5][0] ),
	.OUT(n1326));
   OAI21 U926 (.OUT(n1327),
	.C(n1328),
	.B(n1326),
	.A(n1324));
   AOI21 U927 (.OUT(n1329),
	.C(n1330),
	.B(\mult_20/ab[6][0] ),
	.A(n1327));
   inverter U928 (.IN(\mult_20/ab[7][0] ),
	.OUT(n1331));
   inverter U929 (.IN(\mult_20/ab[4][7] ),
	.OUT(n1332));
   inverter U930 (.IN(\mult_20/ab[5][6] ),
	.OUT(n1333));
   inverter U931 (.IN(\mult_20/ab[5][7] ),
	.OUT(n1334));
   inverter U932 (.IN(\mult_20/ab[6][6] ),
	.OUT(n1335));
   inverter U933 (.IN(\mult_20/ab[7][7] ),
	.OUT(n112));
   AOI21 U934 (.OUT(n1336),
	.C(n1338),
	.B(\mult_20/ab[5][5] ),
	.A(n1337));
   inverter U935 (.IN(\mult_20/ab[6][5] ),
	.OUT(n1339));
   OAI21 U936 (.OUT(n1340),
	.C(n1341),
	.B(n1339),
	.A(n1336));
   AOI21 U937 (.OUT(n1342),
	.C(n1343),
	.B(\mult_20/ab[6][4] ),
	.A(n1297));
   NAND2 U938 (.A(\mult_19_3/ab[0][3] ),
	.B(\mult_19_3/ab[1][2] ),
	.OUT(n1344));
   AOI21 U939 (.OUT(n1345),
	.C(n1347),
	.B(n1346),
	.A(\mult_19_3/ab[2][2] ));
   NAND2 U940 (.A(\mult_19_3/ab[1][3] ),
	.B(\mult_19_3/ab[0][4] ),
	.OUT(n1348));
   inverter U941 (.IN(\mult_19_3/ab[3][2] ),
	.OUT(n1349));
   OAI21 U942 (.OUT(n1350),
	.C(n1351),
	.B(n1349),
	.A(n1345));
   NAND2 U943 (.A(\mult_19_3/ab[1][4] ),
	.B(\mult_19_3/ab[0][5] ),
	.OUT(n1352));
   inverter U944 (.IN(\mult_19_3/ab[3][3] ),
	.OUT(n1353));
   OAI21 U945 (.OUT(n1354),
	.C(n1356),
	.B(n1355),
	.A(n1348));
   AOI21 U946 (.OUT(n1357),
	.C(n1358),
	.B(\mult_19_3/ab[4][2] ),
	.A(n1350));
   NAND2 U947 (.A(\mult_19_3/ab[1][5] ),
	.B(\mult_19_3/ab[0][6] ),
	.OUT(n1359));
   inverter U948 (.IN(\mult_19_3/ab[3][4] ),
	.OUT(n1360));
   OAI21 U949 (.OUT(n1361),
	.C(n1363),
	.B(n1362),
	.A(n1352));
   AOI21 U950 (.OUT(n1364),
	.C(n1365),
	.B(\mult_19_3/ab[3][3] ),
	.A(n1354));
   inverter U951 (.IN(\mult_19_3/ab[5][2] ),
	.OUT(n1366));
   OAI21 U952 (.OUT(n1367),
	.C(n1368),
	.B(n1366),
	.A(n1357));
   NAND2 U953 (.A(\mult_19_3/ab[1][6] ),
	.B(\mult_19_3/ab[0][7] ),
	.OUT(n1369));
   OAI21 U954 (.OUT(n1370),
	.C(n1372),
	.B(n1371),
	.A(n1359));
   inverter U955 (.IN(\mult_19_3/ab[4][4] ),
	.OUT(n1373));
   AOI21 U956 (.OUT(n1374),
	.C(n1375),
	.B(\mult_19_3/ab[3][4] ),
	.A(n1361));
   OAI21 U957 (.OUT(n1376),
	.C(n1378),
	.B(n1377),
	.A(n1364));
   AOI21 U958 (.OUT(n1379),
	.C(n1380),
	.B(\mult_19_3/ab[6][2] ),
	.A(n1367));
   inverter U959 (.IN(\mult_19_3/ab[3][6] ),
	.OUT(n1381));
   inverter U960 (.IN(\mult_19_3/ab[2][7] ),
	.OUT(n1382));
   OAI21 U961 (.OUT(n1383),
	.C(n1386),
	.B(n1385),
	.A(n1384));
   inverter U962 (.IN(\mult_19_3/ab[5][4] ),
	.OUT(n1387));
   AOI21 U963 (.OUT(n1388),
	.C(n1390),
	.B(\mult_19_3/ab[4][4] ),
	.A(n1389));
   AOI21 U964 (.OUT(n1391),
	.C(n1392),
	.B(\mult_19_3/ab[5][3] ),
	.A(n1376));
   inverter U965 (.IN(\mult_19_3/ab[4][6] ),
	.OUT(n1393));
   inverter U966 (.IN(\mult_19_3/ab[3][7] ),
	.OUT(n1394));
   AOI21 U967 (.OUT(n1395),
	.C(n1396),
	.B(\mult_19_3/ab[4][5] ),
	.A(n1383));
   OAI21 U968 (.OUT(n1397),
	.C(n1398),
	.B(n1387),
	.A(n1388));
   OAI21 U969 (.OUT(n1399),
	.C(n1401),
	.B(n1400),
	.A(n1391));
   NAND2 U970 (.A(\mult_19_3/ab[0][2] ),
	.B(\mult_19_3/ab[1][1] ),
	.OUT(n1402));
   OAI21 U971 (.OUT(n1403),
	.C(n1405),
	.B(n1402),
	.A(n1404));
   inverter U972 (.IN(\mult_19_3/ab[3][1] ),
	.OUT(n1406));
   AOI21 U973 (.OUT(n1407),
	.C(n1408),
	.B(\mult_19_3/ab[3][1] ),
	.A(n1403));
   OAI21 U974 (.OUT(n1409),
	.C(n1411),
	.B(n1410),
	.A(n1407));
   AOI21 U975 (.OUT(n1412),
	.C(n1413),
	.B(\mult_19_3/ab[5][1] ),
	.A(n1409));
   inverter U976 (.IN(\mult_19_3/ab[6][1] ),
	.OUT(n1414));
   OAI21 U977 (.OUT(n1415),
	.C(n1416),
	.B(n1414),
	.A(n1412));
   NAND2 U978 (.A(\mult_19_3/ab[0][1] ),
	.B(\mult_19_3/ab[1][0] ),
	.OUT(n1417));
   AOI21 U979 (.OUT(n1418),
	.C(n1420),
	.B(n1419),
	.A(\mult_19_3/ab[2][0] ));
   inverter U980 (.IN(\mult_19_3/ab[3][0] ),
	.OUT(n1421));
   OAI21 U981 (.OUT(n1422),
	.C(n1423),
	.B(n1421),
	.A(n1418));
   AOI21 U982 (.OUT(n1424),
	.C(n1425),
	.B(\mult_19_3/ab[4][0] ),
	.A(n1422));
   inverter U983 (.IN(\mult_19_3/ab[5][0] ),
	.OUT(n1426));
   OAI21 U984 (.OUT(n1427),
	.C(n1428),
	.B(n1426),
	.A(n1424));
   AOI21 U985 (.OUT(n1429),
	.C(n1430),
	.B(\mult_19_3/ab[6][0] ),
	.A(n1427));
   inverter U986 (.IN(\mult_19_3/ab[7][0] ),
	.OUT(n1431));
   inverter U987 (.IN(\mult_19_3/ab[4][7] ),
	.OUT(n1432));
   inverter U988 (.IN(\mult_19_3/ab[5][6] ),
	.OUT(n1433));
   inverter U989 (.IN(\mult_19_3/ab[5][7] ),
	.OUT(n1434));
   inverter U990 (.IN(\mult_19_3/ab[6][6] ),
	.OUT(n1435));
   inverter U991 (.IN(\mult_19_3/ab[7][7] ),
	.OUT(n97));
   AOI21 U992 (.OUT(n1436),
	.C(n1438),
	.B(\mult_19_3/ab[5][5] ),
	.A(n1437));
   inverter U993 (.IN(\mult_19_3/ab[6][5] ),
	.OUT(n1439));
   OAI21 U994 (.OUT(n1440),
	.C(n1441),
	.B(n1439),
	.A(n1436));
   AOI21 U995 (.OUT(n1442),
	.C(n1443),
	.B(\mult_19_3/ab[6][4] ),
	.A(n1397));
   NAND2 U996 (.A(\mult_19_2/ab[0][3] ),
	.B(\mult_19_2/ab[1][2] ),
	.OUT(n1444));
   AOI21 U997 (.OUT(n1445),
	.C(n1447),
	.B(n1446),
	.A(\mult_19_2/ab[2][2] ));
   NAND2 U998 (.A(\mult_19_2/ab[1][3] ),
	.B(\mult_19_2/ab[0][4] ),
	.OUT(n1448));
   inverter U999 (.IN(\mult_19_2/ab[3][2] ),
	.OUT(n1449));
   OAI21 U1000 (.OUT(n1450),
	.C(n1451),
	.B(n1449),
	.A(n1445));
   NAND2 U1001 (.A(\mult_19_2/ab[1][4] ),
	.B(\mult_19_2/ab[0][5] ),
	.OUT(n1452));
   inverter U1002 (.IN(\mult_19_2/ab[3][3] ),
	.OUT(n1453));
   OAI21 U1003 (.OUT(n1454),
	.C(n1456),
	.B(n1455),
	.A(n1448));
   AOI21 U1004 (.OUT(n1457),
	.C(n1458),
	.B(\mult_19_2/ab[4][2] ),
	.A(n1450));
   NAND2 U1005 (.A(\mult_19_2/ab[1][5] ),
	.B(\mult_19_2/ab[0][6] ),
	.OUT(n1459));
   inverter U1006 (.IN(\mult_19_2/ab[3][4] ),
	.OUT(n1460));
   OAI21 U1007 (.OUT(n1461),
	.C(n1463),
	.B(n1462),
	.A(n1452));
   AOI21 U1008 (.OUT(n1464),
	.C(n1465),
	.B(\mult_19_2/ab[3][3] ),
	.A(n1454));
   inverter U1009 (.IN(\mult_19_2/ab[5][2] ),
	.OUT(n1466));
   OAI21 U1010 (.OUT(n1467),
	.C(n1468),
	.B(n1466),
	.A(n1457));
   NAND2 U1011 (.A(\mult_19_2/ab[1][6] ),
	.B(\mult_19_2/ab[0][7] ),
	.OUT(n1469));
   OAI21 U1012 (.OUT(n1470),
	.C(n1472),
	.B(n1471),
	.A(n1459));
   inverter U1013 (.IN(\mult_19_2/ab[4][4] ),
	.OUT(n1473));
   AOI21 U1014 (.OUT(n1474),
	.C(n1475),
	.B(\mult_19_2/ab[3][4] ),
	.A(n1461));
   OAI21 U1015 (.OUT(n1476),
	.C(n1478),
	.B(n1477),
	.A(n1464));
   AOI21 U1016 (.OUT(n1479),
	.C(n1480),
	.B(\mult_19_2/ab[6][2] ),
	.A(n1467));
   inverter U1017 (.IN(\mult_19_2/ab[3][6] ),
	.OUT(n1481));
   inverter U1018 (.IN(\mult_19_2/ab[2][7] ),
	.OUT(n1482));
   OAI21 U1019 (.OUT(n1483),
	.C(n1486),
	.B(n1485),
	.A(n1484));
   inverter U1020 (.IN(\mult_19_2/ab[5][4] ),
	.OUT(n1487));
   AOI21 U1021 (.OUT(n1488),
	.C(n1490),
	.B(\mult_19_2/ab[4][4] ),
	.A(n1489));
   AOI21 U1022 (.OUT(n1491),
	.C(n1492),
	.B(\mult_19_2/ab[5][3] ),
	.A(n1476));
   inverter U1023 (.IN(\mult_19_2/ab[4][6] ),
	.OUT(n1493));
   inverter U1024 (.IN(\mult_19_2/ab[3][7] ),
	.OUT(n1494));
   AOI21 U1025 (.OUT(n1495),
	.C(n1496),
	.B(\mult_19_2/ab[4][5] ),
	.A(n1483));
   OAI21 U1026 (.OUT(n1497),
	.C(n1498),
	.B(n1487),
	.A(n1488));
   OAI21 U1027 (.OUT(n1499),
	.C(n1501),
	.B(n1500),
	.A(n1491));
   NAND2 U1028 (.A(\mult_19_2/ab[0][2] ),
	.B(\mult_19_2/ab[1][1] ),
	.OUT(n1502));
   OAI21 U1029 (.OUT(n1503),
	.C(n1505),
	.B(n1502),
	.A(n1504));
   inverter U1030 (.IN(\mult_19_2/ab[3][1] ),
	.OUT(n1506));
   AOI21 U1031 (.OUT(n1507),
	.C(n1508),
	.B(\mult_19_2/ab[3][1] ),
	.A(n1503));
   OAI21 U1032 (.OUT(n1509),
	.C(n1511),
	.B(n1510),
	.A(n1507));
   AOI21 U1033 (.OUT(n1512),
	.C(n1513),
	.B(\mult_19_2/ab[5][1] ),
	.A(n1509));
   inverter U1034 (.IN(\mult_19_2/ab[6][1] ),
	.OUT(n1514));
   OAI21 U1035 (.OUT(n1515),
	.C(n1516),
	.B(n1514),
	.A(n1512));
   NAND2 U1036 (.A(\mult_19_2/ab[0][1] ),
	.B(\mult_19_2/ab[1][0] ),
	.OUT(n1517));
   AOI21 U1037 (.OUT(n1518),
	.C(n1520),
	.B(n1519),
	.A(\mult_19_2/ab[2][0] ));
   inverter U1038 (.IN(\mult_19_2/ab[3][0] ),
	.OUT(n1521));
   OAI21 U1039 (.OUT(n1522),
	.C(n1523),
	.B(n1521),
	.A(n1518));
   AOI21 U1040 (.OUT(n1524),
	.C(n1525),
	.B(\mult_19_2/ab[4][0] ),
	.A(n1522));
   inverter U1041 (.IN(\mult_19_2/ab[5][0] ),
	.OUT(n1526));
   OAI21 U1042 (.OUT(n1527),
	.C(n1528),
	.B(n1526),
	.A(n1524));
   AOI21 U1043 (.OUT(n1529),
	.C(n1530),
	.B(\mult_19_2/ab[6][0] ),
	.A(n1527));
   inverter U1044 (.IN(\mult_19_2/ab[7][0] ),
	.OUT(n1531));
   inverter U1045 (.IN(\mult_19_2/ab[4][7] ),
	.OUT(n1532));
   inverter U1046 (.IN(\mult_19_2/ab[5][6] ),
	.OUT(n1533));
   inverter U1047 (.IN(\mult_19_2/ab[5][7] ),
	.OUT(n1534));
   inverter U1048 (.IN(\mult_19_2/ab[6][6] ),
	.OUT(n1535));
   inverter U1049 (.IN(\mult_19_2/ab[7][7] ),
	.OUT(n82));
   AOI21 U1050 (.OUT(n1536),
	.C(n1538),
	.B(\mult_19_2/ab[5][5] ),
	.A(n1537));
   inverter U1051 (.IN(\mult_19_2/ab[6][5] ),
	.OUT(n1539));
   OAI21 U1052 (.OUT(n1540),
	.C(n1541),
	.B(n1539),
	.A(n1536));
   AOI21 U1053 (.OUT(n1542),
	.C(n1543),
	.B(\mult_19_2/ab[6][4] ),
	.A(n1497));
   NAND2 U1054 (.A(\mult_19/ab[0][3] ),
	.B(\mult_19/ab[1][2] ),
	.OUT(n1544));
   AOI21 U1055 (.OUT(n1545),
	.C(n1547),
	.B(n1546),
	.A(\mult_19/ab[2][2] ));
   NAND2 U1056 (.A(\mult_19/ab[1][3] ),
	.B(\mult_19/ab[0][4] ),
	.OUT(n1548));
   inverter U1057 (.IN(\mult_19/ab[3][2] ),
	.OUT(n1549));
   OAI21 U1058 (.OUT(n1550),
	.C(n1551),
	.B(n1549),
	.A(n1545));
   NAND2 U1059 (.A(\mult_19/ab[1][4] ),
	.B(\mult_19/ab[0][5] ),
	.OUT(n1552));
   inverter U1060 (.IN(\mult_19/ab[3][3] ),
	.OUT(n1553));
   OAI21 U1061 (.OUT(n1554),
	.C(n1556),
	.B(n1555),
	.A(n1548));
   AOI21 U1062 (.OUT(n1557),
	.C(n1558),
	.B(\mult_19/ab[4][2] ),
	.A(n1550));
   NAND2 U1063 (.A(\mult_19/ab[1][5] ),
	.B(\mult_19/ab[0][6] ),
	.OUT(n1559));
   inverter U1064 (.IN(\mult_19/ab[3][4] ),
	.OUT(n1560));
   OAI21 U1065 (.OUT(n1561),
	.C(n1563),
	.B(n1562),
	.A(n1552));
   AOI21 U1066 (.OUT(n1564),
	.C(n1565),
	.B(\mult_19/ab[3][3] ),
	.A(n1554));
   inverter U1067 (.IN(\mult_19/ab[5][2] ),
	.OUT(n1566));
   OAI21 U1068 (.OUT(n1567),
	.C(n1568),
	.B(n1566),
	.A(n1557));
   NAND2 U1069 (.A(\mult_19/ab[1][6] ),
	.B(\mult_19/ab[0][7] ),
	.OUT(n1569));
   OAI21 U1070 (.OUT(n1570),
	.C(n1572),
	.B(n1571),
	.A(n1559));
   inverter U1071 (.IN(\mult_19/ab[4][4] ),
	.OUT(n1573));
   AOI21 U1072 (.OUT(n1574),
	.C(n1575),
	.B(\mult_19/ab[3][4] ),
	.A(n1561));
   OAI21 U1073 (.OUT(n1576),
	.C(n1578),
	.B(n1577),
	.A(n1564));
   AOI21 U1074 (.OUT(n1579),
	.C(n1580),
	.B(\mult_19/ab[6][2] ),
	.A(n1567));
   inverter U1075 (.IN(\mult_19/ab[3][6] ),
	.OUT(n1581));
   inverter U1076 (.IN(\mult_19/ab[2][7] ),
	.OUT(n1582));
   OAI21 U1077 (.OUT(n1583),
	.C(n1586),
	.B(n1585),
	.A(n1584));
   inverter U1078 (.IN(\mult_19/ab[5][4] ),
	.OUT(n1587));
   AOI21 U1079 (.OUT(n1588),
	.C(n1590),
	.B(\mult_19/ab[4][4] ),
	.A(n1589));
   AOI21 U1080 (.OUT(n1591),
	.C(n1592),
	.B(\mult_19/ab[5][3] ),
	.A(n1576));
   inverter U1081 (.IN(\mult_19/ab[4][6] ),
	.OUT(n1593));
   inverter U1082 (.IN(\mult_19/ab[3][7] ),
	.OUT(n1594));
   AOI21 U1083 (.OUT(n1595),
	.C(n1596),
	.B(\mult_19/ab[4][5] ),
	.A(n1583));
   OAI21 U1084 (.OUT(n1597),
	.C(n1598),
	.B(n1587),
	.A(n1588));
   OAI21 U1085 (.OUT(n1599),
	.C(n1601),
	.B(n1600),
	.A(n1591));
   NAND2 U1086 (.A(\mult_19/ab[0][2] ),
	.B(\mult_19/ab[1][1] ),
	.OUT(n1602));
   OAI21 U1087 (.OUT(n1603),
	.C(n1605),
	.B(n1602),
	.A(n1604));
   inverter U1088 (.IN(\mult_19/ab[3][1] ),
	.OUT(n1606));
   AOI21 U1089 (.OUT(n1607),
	.C(n1608),
	.B(\mult_19/ab[3][1] ),
	.A(n1603));
   OAI21 U1090 (.OUT(n1609),
	.C(n1611),
	.B(n1610),
	.A(n1607));
   AOI21 U1091 (.OUT(n1612),
	.C(n1613),
	.B(\mult_19/ab[5][1] ),
	.A(n1609));
   inverter U1092 (.IN(\mult_19/ab[6][1] ),
	.OUT(n1614));
   OAI21 U1093 (.OUT(n1615),
	.C(n1616),
	.B(n1614),
	.A(n1612));
   NAND2 U1094 (.A(\mult_19/ab[0][1] ),
	.B(\mult_19/ab[1][0] ),
	.OUT(n1617));
   AOI21 U1095 (.OUT(n1618),
	.C(n1620),
	.B(n1619),
	.A(\mult_19/ab[2][0] ));
   inverter U1096 (.IN(\mult_19/ab[3][0] ),
	.OUT(n1621));
   OAI21 U1097 (.OUT(n1622),
	.C(n1623),
	.B(n1621),
	.A(n1618));
   AOI21 U1098 (.OUT(n1624),
	.C(n1625),
	.B(\mult_19/ab[4][0] ),
	.A(n1622));
   inverter U1099 (.IN(\mult_19/ab[5][0] ),
	.OUT(n1626));
   OAI21 U1100 (.OUT(n1627),
	.C(n1628),
	.B(n1626),
	.A(n1624));
   AOI21 U1101 (.OUT(n1629),
	.C(n1630),
	.B(\mult_19/ab[6][0] ),
	.A(n1627));
   inverter U1102 (.IN(\mult_19/ab[7][0] ),
	.OUT(n1631));
   inverter U1103 (.IN(\mult_19/ab[4][7] ),
	.OUT(n1632));
   inverter U1104 (.IN(\mult_19/ab[5][6] ),
	.OUT(n1633));
   inverter U1105 (.IN(\mult_19/ab[5][7] ),
	.OUT(n1634));
   inverter U1106 (.IN(\mult_19/ab[6][6] ),
	.OUT(n1635));
   inverter U1107 (.IN(\mult_19/ab[7][7] ),
	.OUT(n67));
   AOI21 U1108 (.OUT(n1636),
	.C(n1638),
	.B(\mult_19/ab[5][5] ),
	.A(n1637));
   inverter U1109 (.IN(\mult_19/ab[6][5] ),
	.OUT(n1639));
   OAI21 U1110 (.OUT(n1640),
	.C(n1641),
	.B(n1639),
	.A(n1636));
   AOI21 U1111 (.OUT(n1642),
	.C(n1643),
	.B(\mult_19/ab[6][4] ),
	.A(n1597));
   NAND2 U1112 (.A(N1),
	.B(N17),
	.OUT(n1644));
   NAND2 U1113 (.A(N49),
	.B(n728),
	.OUT(n1645));
   OAI21 U1114 (.OUT(n1646),
	.C(n1648),
	.B(n1645),
	.A(n1647));
   AOI21 U1115 (.OUT(n1649),
	.C(n1650),
	.B(N51),
	.A(n1646));
   inverter U1116 (.IN(N52),
	.OUT(n1651));
   OAI21 U1117 (.OUT(n1652),
	.C(n1653),
	.B(n1651),
	.A(n1649));
   inverter U1118 (.IN(N53),
	.OUT(n1654));
   AOI21 U1119 (.OUT(n1655),
	.C(n1656),
	.B(N53),
	.A(n1652));
   inverter U1120 (.IN(N54),
	.OUT(n1657));
   AOI21 U1121 (.OUT(n1658),
	.C(n1660),
	.B(N54),
	.A(n1659));
   inverter U1122 (.IN(N55),
	.OUT(n1661));
   AOI21 U1123 (.OUT(n1662),
	.C(n1664),
	.B(N55),
	.A(n1663));
   inverter U1124 (.IN(N56),
	.OUT(n1665));
   AOI21 U1125 (.OUT(n1666),
	.C(n1668),
	.B(N56),
	.A(n1667));
   inverter U1126 (.IN(N57),
	.OUT(n1669));
   AOI21 U1127 (.OUT(n1670),
	.C(n1672),
	.B(N57),
	.A(n1671));
   inverter U1128 (.IN(N58),
	.OUT(n1673));
   AOI21 U1129 (.OUT(n1674),
	.C(n1676),
	.B(N58),
	.A(n1675));
   inverter U1130 (.IN(N59),
	.OUT(n1677));
   AOI21 U1131 (.OUT(n1678),
	.C(n1680),
	.B(N59),
	.A(n1679));
   inverter U1132 (.IN(N60),
	.OUT(n1681));
   AOI21 U1133 (.OUT(n1682),
	.C(n1684),
	.B(N60),
	.A(n1683));
   inverter U1134 (.IN(N61),
	.OUT(n1685));
   AOI21 U1135 (.OUT(n1686),
	.C(n1688),
	.B(N61),
	.A(n1687));
   inverter U1136 (.IN(N62),
	.OUT(n1689));
   AOI21 U1137 (.OUT(n206),
	.C(n1691),
	.B(N62),
	.A(n1690));
   inverter U1138 (.IN(N63),
	.OUT(n207));
   NAND2 U1139 (.A(N161),
	.B(N177),
	.OUT(n1692));
   NAND2 U1140 (.A(N209),
	.B(n734),
	.OUT(n1693));
   OAI21 U1141 (.OUT(n1694),
	.C(n1696),
	.B(n1693),
	.A(n1695));
   AOI21 U1142 (.OUT(n1697),
	.C(n1698),
	.B(N211),
	.A(n1694));
   inverter U1143 (.IN(N212),
	.OUT(n1699));
   OAI21 U1144 (.OUT(n1700),
	.C(n1701),
	.B(n1699),
	.A(n1697));
   inverter U1145 (.IN(N213),
	.OUT(n1702));
   AOI21 U1146 (.OUT(n1703),
	.C(n1704),
	.B(N213),
	.A(n1700));
   inverter U1147 (.IN(N214),
	.OUT(n1705));
   AOI21 U1148 (.OUT(n1706),
	.C(n1708),
	.B(N214),
	.A(n1707));
   inverter U1149 (.IN(N215),
	.OUT(n1709));
   AOI21 U1150 (.OUT(n1710),
	.C(n1712),
	.B(N215),
	.A(n1711));
   inverter U1151 (.IN(N216),
	.OUT(n1713));
   AOI21 U1152 (.OUT(n1714),
	.C(n1716),
	.B(N216),
	.A(n1715));
   inverter U1153 (.IN(N217),
	.OUT(n1717));
   AOI21 U1154 (.OUT(n1718),
	.C(n1720),
	.B(N217),
	.A(n1719));
   inverter U1155 (.IN(N218),
	.OUT(n1721));
   AOI21 U1156 (.OUT(n1722),
	.C(n1724),
	.B(N218),
	.A(n1723));
   inverter U1157 (.IN(N219),
	.OUT(n1725));
   AOI21 U1158 (.OUT(n1726),
	.C(n1728),
	.B(N219),
	.A(n1727));
   inverter U1159 (.IN(N220),
	.OUT(n1729));
   AOI21 U1160 (.OUT(n1730),
	.C(n1732),
	.B(N220),
	.A(n1731));
   inverter U1161 (.IN(N221),
	.OUT(n1733));
   AOI21 U1162 (.OUT(n1734),
	.C(n1736),
	.B(N221),
	.A(n1735));
   inverter U1163 (.IN(N222),
	.OUT(n1737));
   AOI21 U1164 (.OUT(n216),
	.C(n1739),
	.B(N222),
	.A(n1738));
   inverter U1165 (.IN(N223),
	.OUT(n217));
   NAND2 U1166 (.A(N81),
	.B(N97),
	.OUT(n1740));
   NAND2 U1167 (.A(N129),
	.B(n740),
	.OUT(n1741));
   OAI21 U1168 (.OUT(n1742),
	.C(n1744),
	.B(n1741),
	.A(n1743));
   AOI21 U1169 (.OUT(n1745),
	.C(n1746),
	.B(N131),
	.A(n1742));
   inverter U1170 (.IN(N132),
	.OUT(n1747));
   OAI21 U1171 (.OUT(n1748),
	.C(n1749),
	.B(n1747),
	.A(n1745));
   inverter U1172 (.IN(N133),
	.OUT(n1750));
   AOI21 U1173 (.OUT(n1751),
	.C(n1752),
	.B(N133),
	.A(n1748));
   inverter U1174 (.IN(N134),
	.OUT(n1753));
   AOI21 U1175 (.OUT(n1754),
	.C(n1756),
	.B(N134),
	.A(n1755));
   inverter U1176 (.IN(N135),
	.OUT(n1757));
   AOI21 U1177 (.OUT(n1758),
	.C(n1760),
	.B(N135),
	.A(n1759));
   inverter U1178 (.IN(N136),
	.OUT(n1761));
   AOI21 U1179 (.OUT(n1762),
	.C(n1764),
	.B(N136),
	.A(n1763));
   inverter U1180 (.IN(N137),
	.OUT(n1765));
   AOI21 U1181 (.OUT(n1766),
	.C(n1768),
	.B(N137),
	.A(n1767));
   inverter U1182 (.IN(N138),
	.OUT(n1769));
   AOI21 U1183 (.OUT(n1770),
	.C(n1772),
	.B(N138),
	.A(n1771));
   inverter U1184 (.IN(N139),
	.OUT(n1773));
   AOI21 U1185 (.OUT(n1774),
	.C(n1776),
	.B(N139),
	.A(n1775));
   inverter U1186 (.IN(N140),
	.OUT(n1777));
   AOI21 U1187 (.OUT(n1778),
	.C(n1780),
	.B(N140),
	.A(n1779));
   inverter U1188 (.IN(N141),
	.OUT(n1781));
   AOI21 U1189 (.OUT(n1782),
	.C(n1784),
	.B(N141),
	.A(n1783));
   inverter U1190 (.IN(N142),
	.OUT(n1785));
   AOI21 U1191 (.OUT(n226),
	.C(n1787),
	.B(N142),
	.A(n1786));
   inverter U1192 (.IN(N143),
	.OUT(n227));
   XOR2 U1193 (.A(n193),
	.B(n194),
	.OUT(\mult_21_3/A1[9] ));
   XOR2 U1194 (.A(n197),
	.B(n198),
	.OUT(\mult_21_3/A1[7] ));
   XOR2 U1195 (.A(n199),
	.B(n200),
	.OUT(\mult_21_3/A1[6] ));
   XOR2 U1196 (.A(n1788),
	.B(n1789),
	.OUT(\mult_21_3/A1[4] ));
   XOR2 U1197 (.A(n1790),
	.B(n1791),
	.OUT(\mult_21_3/A1[2] ));
   XOR2 U1198 (.A(n188),
	.B(n189),
	.OUT(\mult_21_3/A1[11] ));
   XOR2 U1199 (.A(n269),
	.B(n1792),
	.OUT(\mult_21_3/A1[0] ));
   XOR2 U1200 (.A(n178),
	.B(n179),
	.OUT(\mult_21_2/A1[9] ));
   XOR2 U1201 (.A(n182),
	.B(n183),
	.OUT(\mult_21_2/A1[7] ));
   XOR2 U1202 (.A(n184),
	.B(n185),
	.OUT(\mult_21_2/A1[6] ));
   XOR2 U1203 (.A(n1793),
	.B(n1794),
	.OUT(\mult_21_2/A1[4] ));
   XOR2 U1204 (.A(n1795),
	.B(n1796),
	.OUT(\mult_21_2/A1[2] ));
   XOR2 U1205 (.A(n173),
	.B(n174),
	.OUT(\mult_21_2/A1[11] ));
   XOR2 U1206 (.A(n324),
	.B(n1797),
	.OUT(\mult_21_2/A1[0] ));
   XOR2 U1207 (.A(n163),
	.B(n164),
	.OUT(\mult_21/A1[9] ));
   XOR2 U1208 (.A(n167),
	.B(n168),
	.OUT(\mult_21/A1[7] ));
   XOR2 U1209 (.A(n169),
	.B(n170),
	.OUT(\mult_21/A1[6] ));
   XOR2 U1210 (.A(n1798),
	.B(n1799),
	.OUT(\mult_21/A1[4] ));
   XOR2 U1211 (.A(n1800),
	.B(n1801),
	.OUT(\mult_21/A1[2] ));
   XOR2 U1212 (.A(n158),
	.B(n159),
	.OUT(\mult_21/A1[11] ));
   XOR2 U1213 (.A(n379),
	.B(n1802),
	.OUT(\mult_21/A1[0] ));
   XOR2 U1214 (.A(n148),
	.B(n149),
	.OUT(\mult_20_3/A1[9] ));
   XOR2 U1215 (.A(n152),
	.B(n153),
	.OUT(\mult_20_3/A1[7] ));
   XOR2 U1216 (.A(n154),
	.B(n155),
	.OUT(\mult_20_3/A1[6] ));
   XOR2 U1217 (.A(n1803),
	.B(n1804),
	.OUT(\mult_20_3/A1[4] ));
   XOR2 U1218 (.A(n1805),
	.B(n1806),
	.OUT(\mult_20_3/A1[2] ));
   XOR2 U1219 (.A(n143),
	.B(n144),
	.OUT(\mult_20_3/A1[11] ));
   XOR2 U1220 (.A(n434),
	.B(n1807),
	.OUT(\mult_20_3/A1[0] ));
   XOR2 U1221 (.A(n133),
	.B(n134),
	.OUT(\mult_20_2/A1[9] ));
   XOR2 U1222 (.A(n137),
	.B(n138),
	.OUT(\mult_20_2/A1[7] ));
   XOR2 U1223 (.A(n139),
	.B(n140),
	.OUT(\mult_20_2/A1[6] ));
   XOR2 U1224 (.A(n1808),
	.B(n1809),
	.OUT(\mult_20_2/A1[4] ));
   XOR2 U1225 (.A(n1810),
	.B(n1811),
	.OUT(\mult_20_2/A1[2] ));
   XOR2 U1226 (.A(n128),
	.B(n129),
	.OUT(\mult_20_2/A1[11] ));
   XOR2 U1227 (.A(n489),
	.B(n1812),
	.OUT(\mult_20_2/A1[0] ));
   XOR2 U1228 (.A(n118),
	.B(n119),
	.OUT(\mult_20/A1[9] ));
   XOR2 U1229 (.A(n122),
	.B(n123),
	.OUT(\mult_20/A1[7] ));
   XOR2 U1230 (.A(n124),
	.B(n125),
	.OUT(\mult_20/A1[6] ));
   XOR2 U1231 (.A(n1813),
	.B(n1814),
	.OUT(\mult_20/A1[4] ));
   XOR2 U1232 (.A(n1815),
	.B(n1816),
	.OUT(\mult_20/A1[2] ));
   XOR2 U1233 (.A(n113),
	.B(n114),
	.OUT(\mult_20/A1[11] ));
   XOR2 U1234 (.A(n544),
	.B(n1817),
	.OUT(\mult_20/A1[0] ));
   XOR2 U1235 (.A(n103),
	.B(n104),
	.OUT(\mult_19_3/A1[9] ));
   XOR2 U1236 (.A(n107),
	.B(n108),
	.OUT(\mult_19_3/A1[7] ));
   XOR2 U1237 (.A(n109),
	.B(n110),
	.OUT(\mult_19_3/A1[6] ));
   XOR2 U1238 (.A(n1818),
	.B(n1819),
	.OUT(\mult_19_3/A1[4] ));
   XOR2 U1239 (.A(n1820),
	.B(n1821),
	.OUT(\mult_19_3/A1[2] ));
   XOR2 U1240 (.A(n98),
	.B(n99),
	.OUT(\mult_19_3/A1[11] ));
   XOR2 U1241 (.A(n599),
	.B(n1822),
	.OUT(\mult_19_3/A1[0] ));
   XOR2 U1242 (.A(n88),
	.B(n89),
	.OUT(\mult_19_2/A1[9] ));
   XOR2 U1243 (.A(n92),
	.B(n93),
	.OUT(\mult_19_2/A1[7] ));
   XOR2 U1244 (.A(n94),
	.B(n95),
	.OUT(\mult_19_2/A1[6] ));
   XOR2 U1245 (.A(n1823),
	.B(n1824),
	.OUT(\mult_19_2/A1[4] ));
   XOR2 U1246 (.A(n1825),
	.B(n1826),
	.OUT(\mult_19_2/A1[2] ));
   XOR2 U1247 (.A(n83),
	.B(n84),
	.OUT(\mult_19_2/A1[11] ));
   XOR2 U1248 (.A(n654),
	.B(n1827),
	.OUT(\mult_19_2/A1[0] ));
   XOR2 U1249 (.A(n73),
	.B(n74),
	.OUT(\mult_19/A1[9] ));
   XOR2 U1250 (.A(n77),
	.B(n78),
	.OUT(\mult_19/A1[7] ));
   XOR2 U1251 (.A(n79),
	.B(n80),
	.OUT(\mult_19/A1[6] ));
   XOR2 U1252 (.A(n1828),
	.B(n1829),
	.OUT(\mult_19/A1[4] ));
   XOR2 U1253 (.A(n1830),
	.B(n1831),
	.OUT(\mult_19/A1[2] ));
   XOR2 U1254 (.A(n68),
	.B(n69),
	.OUT(\mult_19/A1[11] ));
   XOR2 U1255 (.A(n709),
	.B(n1832),
	.OUT(\mult_19/A1[0] ));
   XOR2 U1256 (.A(n1833),
	.B(n1834),
	.OUT(N80));
   XOR2 U1257 (.A(n208),
	.B(n1835),
	.OUT(N79));
   XOR2 U1258 (.A(n1836),
	.B(n1837),
	.OUT(N78));
   XOR2 U1259 (.A(n1838),
	.B(n1839),
	.OUT(N77));
   XOR2 U1260 (.A(n1840),
	.B(n1841),
	.OUT(N76));
   XOR2 U1261 (.A(n1842),
	.B(n1843),
	.OUT(N75));
   XOR2 U1262 (.A(n1844),
	.B(n1845),
	.OUT(N74));
   XOR2 U1263 (.A(n1846),
	.B(n1847),
	.OUT(N73));
   XOR2 U1264 (.A(n1848),
	.B(n1849),
	.OUT(N72));
   XOR2 U1265 (.A(n1850),
	.B(n1851),
	.OUT(N71));
   XOR2 U1266 (.A(n1852),
	.B(n1853),
	.OUT(N70));
   XOR2 U1267 (.A(n1854),
	.B(n1855),
	.OUT(N69));
   XOR2 U1268 (.A(n1856),
	.B(n1857),
	.OUT(N68));
   XOR2 U1269 (.A(n1858),
	.B(n1859),
	.OUT(N67));
   XOR2 U1270 (.A(n730),
	.B(n1860),
	.OUT(N66));
   XOR2 U1271 (.A(N49),
	.B(n728),
	.OUT(N65));
   XOR2 U1272 (.A(n1861),
	.B(n1862),
	.OUT(N240));
   XOR2 U1273 (.A(n218),
	.B(n1863),
	.OUT(N239));
   XOR2 U1274 (.A(n1864),
	.B(n1865),
	.OUT(N238));
   XOR2 U1275 (.A(n1866),
	.B(n1867),
	.OUT(N237));
   XOR2 U1276 (.A(n1868),
	.B(n1869),
	.OUT(N236));
   XOR2 U1277 (.A(n1870),
	.B(n1871),
	.OUT(N235));
   XOR2 U1278 (.A(n1872),
	.B(n1873),
	.OUT(N234));
   XOR2 U1279 (.A(n1874),
	.B(n1875),
	.OUT(N233));
   XOR2 U1280 (.A(n1876),
	.B(n1877),
	.OUT(N232));
   XOR2 U1281 (.A(n1878),
	.B(n1879),
	.OUT(N231));
   XOR2 U1282 (.A(n1880),
	.B(n1881),
	.OUT(N230));
   XOR2 U1283 (.A(n1882),
	.B(n1883),
	.OUT(N229));
   XOR2 U1284 (.A(n1884),
	.B(n1885),
	.OUT(N228));
   XOR2 U1285 (.A(n1886),
	.B(n1887),
	.OUT(N227));
   XOR2 U1286 (.A(n736),
	.B(n1888),
	.OUT(N226));
   XOR2 U1287 (.A(N209),
	.B(n734),
	.OUT(N225));
   XOR2 U1288 (.A(n1889),
	.B(n1890),
	.OUT(N160));
   XOR2 U1289 (.A(n228),
	.B(n1891),
	.OUT(N159));
   XOR2 U1290 (.A(n1892),
	.B(n1893),
	.OUT(N158));
   XOR2 U1291 (.A(n1894),
	.B(n1895),
	.OUT(N157));
   XOR2 U1292 (.A(n1896),
	.B(n1897),
	.OUT(N156));
   XOR2 U1293 (.A(n1898),
	.B(n1899),
	.OUT(N155));
   XOR2 U1294 (.A(n1900),
	.B(n1901),
	.OUT(N154));
   XOR2 U1295 (.A(n1902),
	.B(n1903),
	.OUT(N153));
   XOR2 U1296 (.A(n1904),
	.B(n1905),
	.OUT(N152));
   XOR2 U1297 (.A(n1906),
	.B(n1907),
	.OUT(N151));
   XOR2 U1298 (.A(n1908),
	.B(n1909),
	.OUT(N150));
   XOR2 U1299 (.A(n1910),
	.B(n1911),
	.OUT(N149));
   XOR2 U1300 (.A(n1912),
	.B(n1913),
	.OUT(N148));
   XOR2 U1301 (.A(n1914),
	.B(n1915),
	.OUT(N147));
   XOR2 U1302 (.A(n742),
	.B(n1916),
	.OUT(N146));
   XOR2 U1303 (.A(N129),
	.B(n740),
	.OUT(N145));
   XOR2 U1304 (.A(n753),
	.B(n754),
	.OUT(n1917));
   XOR2 U1305 (.A(n760),
	.B(n761),
	.OUT(n1918));
   XOR2 U1306 (.A(n777),
	.B(n1919),
	.OUT(n248));
   XOR2 U1307 (.A(n1920),
	.B(\mult_21_3/ab[2][6] ),
	.OUT(n232));
   XOR2 U1308 (.A(n785),
	.B(n770),
	.OUT(n1921));
   XOR2 U1309 (.A(\mult_21_3/ab[4][4] ),
	.B(n774),
	.OUT(n239));
   XOR2 U1310 (.A(\mult_21_3/ab[5][3] ),
	.B(n776),
	.OUT(n1922));
   XOR2 U1311 (.A(\mult_21_3/ab[4][5] ),
	.B(n783),
	.OUT(n251));
   XOR2 U1312 (.A(\mult_21_3/ab[5][4] ),
	.B(n788),
	.OUT(n1923));
   XOR2 U1313 (.A(\mult_21_3/ab[6][3] ),
	.B(n791),
	.OUT(n254));
   XOR2 U1314 (.A(n1924),
	.B(n837),
	.OUT(n257));
   XOR2 U1315 (.A(\mult_21_3/ab[6][4] ),
	.B(n797),
	.OUT(n1925));
   XOR2 U1316 (.A(\mult_21_3/ab[7][3] ),
	.B(n799),
	.OUT(n259));
   XOR2 U1317 (.A(\mult_21_3/ab[3][2] ),
	.B(n745),
	.OUT(n1926));
   XOR2 U1318 (.A(\mult_21_3/ab[4][2] ),
	.B(n750),
	.OUT(n265));
   XOR2 U1319 (.A(\mult_21_3/ab[5][2] ),
	.B(n757),
	.OUT(n1927));
   XOR2 U1320 (.A(\mult_21_3/ab[6][2] ),
	.B(n767),
	.OUT(n268));
   XOR2 U1321 (.A(\mult_21_3/ab[7][2] ),
	.B(n779),
	.OUT(n1928));
   XOR2 U1322 (.A(n806),
	.B(n803),
	.OUT(n1929));
   XOR2 U1323 (.A(\mult_21_3/ab[4][1] ),
	.B(n807),
	.OUT(n274));
   XOR2 U1324 (.A(\mult_21_3/ab[5][1] ),
	.B(n809),
	.OUT(n1930));
   XOR2 U1325 (.A(\mult_21_3/ab[6][1] ),
	.B(n812),
	.OUT(n277));
   XOR2 U1326 (.A(\mult_21_3/ab[7][1] ),
	.B(n815),
	.OUT(n1931));
   XOR2 U1327 (.A(\mult_21_3/ab[6][5] ),
	.B(n836),
	.OUT(n280));
   XOR2 U1328 (.A(\mult_21_3/ab[7][5] ),
	.B(n840),
	.OUT(n282));
   XOR2 U1329 (.A(\mult_21_3/ab[7][4] ),
	.B(n842),
	.OUT(n1932));
   XOR2 U1330 (.A(\mult_21_3/ab[7][0] ),
	.B(n829),
	.OUT(n283));
   XOR2 U1331 (.A(\mult_21_3/ab[6][0] ),
	.B(n827),
	.OUT(n1789));
   XOR2 U1332 (.A(\mult_21_3/ab[5][0] ),
	.B(n824),
	.OUT(n284));
   XOR2 U1333 (.A(\mult_21_3/ab[4][0] ),
	.B(n822),
	.OUT(n1791));
   XOR2 U1334 (.A(\mult_21_3/ab[3][0] ),
	.B(n818),
	.OUT(n285));
   XOR2 U1335 (.A(n819),
	.B(\mult_21_3/ab[2][0] ),
	.OUT(n1792));
   XOR2 U1336 (.A(n853),
	.B(n854),
	.OUT(n1933));
   XOR2 U1337 (.A(n860),
	.B(n861),
	.OUT(n1934));
   XOR2 U1338 (.A(n877),
	.B(n1935),
	.OUT(n303));
   XOR2 U1339 (.A(n1936),
	.B(\mult_21_2/ab[2][6] ),
	.OUT(n287));
   XOR2 U1340 (.A(n885),
	.B(n870),
	.OUT(n1937));
   XOR2 U1341 (.A(\mult_21_2/ab[4][4] ),
	.B(n874),
	.OUT(n294));
   XOR2 U1342 (.A(\mult_21_2/ab[5][3] ),
	.B(n876),
	.OUT(n1938));
   XOR2 U1343 (.A(\mult_21_2/ab[4][5] ),
	.B(n883),
	.OUT(n306));
   XOR2 U1344 (.A(\mult_21_2/ab[5][4] ),
	.B(n888),
	.OUT(n1939));
   XOR2 U1345 (.A(\mult_21_2/ab[6][3] ),
	.B(n891),
	.OUT(n309));
   XOR2 U1346 (.A(n1940),
	.B(n937),
	.OUT(n312));
   XOR2 U1347 (.A(\mult_21_2/ab[6][4] ),
	.B(n897),
	.OUT(n1941));
   XOR2 U1348 (.A(\mult_21_2/ab[7][3] ),
	.B(n899),
	.OUT(n314));
   XOR2 U1349 (.A(\mult_21_2/ab[3][2] ),
	.B(n845),
	.OUT(n1942));
   XOR2 U1350 (.A(\mult_21_2/ab[4][2] ),
	.B(n850),
	.OUT(n320));
   XOR2 U1351 (.A(\mult_21_2/ab[5][2] ),
	.B(n857),
	.OUT(n1943));
   XOR2 U1352 (.A(\mult_21_2/ab[6][2] ),
	.B(n867),
	.OUT(n323));
   XOR2 U1353 (.A(\mult_21_2/ab[7][2] ),
	.B(n879),
	.OUT(n1944));
   XOR2 U1354 (.A(n906),
	.B(n903),
	.OUT(n1945));
   XOR2 U1355 (.A(\mult_21_2/ab[4][1] ),
	.B(n907),
	.OUT(n329));
   XOR2 U1356 (.A(\mult_21_2/ab[5][1] ),
	.B(n909),
	.OUT(n1946));
   XOR2 U1357 (.A(\mult_21_2/ab[6][1] ),
	.B(n912),
	.OUT(n332));
   XOR2 U1358 (.A(\mult_21_2/ab[7][1] ),
	.B(n915),
	.OUT(n1947));
   XOR2 U1359 (.A(\mult_21_2/ab[6][5] ),
	.B(n936),
	.OUT(n335));
   XOR2 U1360 (.A(\mult_21_2/ab[7][5] ),
	.B(n940),
	.OUT(n337));
   XOR2 U1361 (.A(\mult_21_2/ab[7][4] ),
	.B(n942),
	.OUT(n1948));
   XOR2 U1362 (.A(\mult_21_2/ab[7][0] ),
	.B(n929),
	.OUT(n338));
   XOR2 U1363 (.A(\mult_21_2/ab[6][0] ),
	.B(n927),
	.OUT(n1794));
   XOR2 U1364 (.A(\mult_21_2/ab[5][0] ),
	.B(n924),
	.OUT(n339));
   XOR2 U1365 (.A(\mult_21_2/ab[4][0] ),
	.B(n922),
	.OUT(n1796));
   XOR2 U1366 (.A(\mult_21_2/ab[3][0] ),
	.B(n918),
	.OUT(n340));
   XOR2 U1367 (.A(n919),
	.B(\mult_21_2/ab[2][0] ),
	.OUT(n1797));
   XOR2 U1368 (.A(n953),
	.B(n954),
	.OUT(n1949));
   XOR2 U1369 (.A(n960),
	.B(n961),
	.OUT(n1950));
   XOR2 U1370 (.A(n977),
	.B(n1951),
	.OUT(n358));
   XOR2 U1371 (.A(n1952),
	.B(\mult_21/ab[2][6] ),
	.OUT(n342));
   XOR2 U1372 (.A(n985),
	.B(n970),
	.OUT(n1953));
   XOR2 U1373 (.A(\mult_21/ab[4][4] ),
	.B(n974),
	.OUT(n349));
   XOR2 U1374 (.A(\mult_21/ab[5][3] ),
	.B(n976),
	.OUT(n1954));
   XOR2 U1375 (.A(\mult_21/ab[4][5] ),
	.B(n983),
	.OUT(n361));
   XOR2 U1376 (.A(\mult_21/ab[5][4] ),
	.B(n988),
	.OUT(n1955));
   XOR2 U1377 (.A(\mult_21/ab[6][3] ),
	.B(n991),
	.OUT(n364));
   XOR2 U1378 (.A(n1956),
	.B(n1037),
	.OUT(n367));
   XOR2 U1379 (.A(\mult_21/ab[6][4] ),
	.B(n997),
	.OUT(n1957));
   XOR2 U1380 (.A(\mult_21/ab[7][3] ),
	.B(n999),
	.OUT(n369));
   XOR2 U1381 (.A(\mult_21/ab[3][2] ),
	.B(n945),
	.OUT(n1958));
   XOR2 U1382 (.A(\mult_21/ab[4][2] ),
	.B(n950),
	.OUT(n375));
   XOR2 U1383 (.A(\mult_21/ab[5][2] ),
	.B(n957),
	.OUT(n1959));
   XOR2 U1384 (.A(\mult_21/ab[6][2] ),
	.B(n967),
	.OUT(n378));
   XOR2 U1385 (.A(\mult_21/ab[7][2] ),
	.B(n979),
	.OUT(n1960));
   XOR2 U1386 (.A(n1006),
	.B(n1003),
	.OUT(n1961));
   XOR2 U1387 (.A(\mult_21/ab[4][1] ),
	.B(n1007),
	.OUT(n384));
   XOR2 U1388 (.A(\mult_21/ab[5][1] ),
	.B(n1009),
	.OUT(n1962));
   XOR2 U1389 (.A(\mult_21/ab[6][1] ),
	.B(n1012),
	.OUT(n387));
   XOR2 U1390 (.A(\mult_21/ab[7][1] ),
	.B(n1015),
	.OUT(n1963));
   XOR2 U1391 (.A(\mult_21/ab[6][5] ),
	.B(n1036),
	.OUT(n390));
   XOR2 U1392 (.A(\mult_21/ab[7][5] ),
	.B(n1040),
	.OUT(n392));
   XOR2 U1393 (.A(\mult_21/ab[7][4] ),
	.B(n1042),
	.OUT(n1964));
   XOR2 U1394 (.A(\mult_21/ab[7][0] ),
	.B(n1029),
	.OUT(n393));
   XOR2 U1395 (.A(\mult_21/ab[6][0] ),
	.B(n1027),
	.OUT(n1799));
   XOR2 U1396 (.A(\mult_21/ab[5][0] ),
	.B(n1024),
	.OUT(n394));
   XOR2 U1397 (.A(\mult_21/ab[4][0] ),
	.B(n1022),
	.OUT(n1801));
   XOR2 U1398 (.A(\mult_21/ab[3][0] ),
	.B(n1018),
	.OUT(n395));
   XOR2 U1399 (.A(n1019),
	.B(\mult_21/ab[2][0] ),
	.OUT(n1802));
   XOR2 U1400 (.A(n1053),
	.B(n1054),
	.OUT(n1965));
   XOR2 U1401 (.A(n1060),
	.B(n1061),
	.OUT(n1966));
   XOR2 U1402 (.A(n1077),
	.B(n1967),
	.OUT(n413));
   XOR2 U1403 (.A(n1968),
	.B(\mult_20_3/ab[2][6] ),
	.OUT(n397));
   XOR2 U1404 (.A(n1085),
	.B(n1070),
	.OUT(n1969));
   XOR2 U1405 (.A(\mult_20_3/ab[4][4] ),
	.B(n1074),
	.OUT(n404));
   XOR2 U1406 (.A(\mult_20_3/ab[5][3] ),
	.B(n1076),
	.OUT(n1970));
   XOR2 U1407 (.A(\mult_20_3/ab[4][5] ),
	.B(n1083),
	.OUT(n416));
   XOR2 U1408 (.A(\mult_20_3/ab[5][4] ),
	.B(n1088),
	.OUT(n1971));
   XOR2 U1409 (.A(\mult_20_3/ab[6][3] ),
	.B(n1091),
	.OUT(n419));
   XOR2 U1410 (.A(n1972),
	.B(n1137),
	.OUT(n422));
   XOR2 U1411 (.A(\mult_20_3/ab[6][4] ),
	.B(n1097),
	.OUT(n1973));
   XOR2 U1412 (.A(\mult_20_3/ab[7][3] ),
	.B(n1099),
	.OUT(n424));
   XOR2 U1413 (.A(\mult_20_3/ab[3][2] ),
	.B(n1045),
	.OUT(n1974));
   XOR2 U1414 (.A(\mult_20_3/ab[4][2] ),
	.B(n1050),
	.OUT(n430));
   XOR2 U1415 (.A(\mult_20_3/ab[5][2] ),
	.B(n1057),
	.OUT(n1975));
   XOR2 U1416 (.A(\mult_20_3/ab[6][2] ),
	.B(n1067),
	.OUT(n433));
   XOR2 U1417 (.A(\mult_20_3/ab[7][2] ),
	.B(n1079),
	.OUT(n1976));
   XOR2 U1418 (.A(n1106),
	.B(n1103),
	.OUT(n1977));
   XOR2 U1419 (.A(\mult_20_3/ab[4][1] ),
	.B(n1107),
	.OUT(n439));
   XOR2 U1420 (.A(\mult_20_3/ab[5][1] ),
	.B(n1109),
	.OUT(n1978));
   XOR2 U1421 (.A(\mult_20_3/ab[6][1] ),
	.B(n1112),
	.OUT(n442));
   XOR2 U1422 (.A(\mult_20_3/ab[7][1] ),
	.B(n1115),
	.OUT(n1979));
   XOR2 U1423 (.A(\mult_20_3/ab[6][5] ),
	.B(n1136),
	.OUT(n445));
   XOR2 U1424 (.A(\mult_20_3/ab[7][5] ),
	.B(n1140),
	.OUT(n447));
   XOR2 U1425 (.A(\mult_20_3/ab[7][4] ),
	.B(n1142),
	.OUT(n1980));
   XOR2 U1426 (.A(\mult_20_3/ab[7][0] ),
	.B(n1129),
	.OUT(n448));
   XOR2 U1427 (.A(\mult_20_3/ab[6][0] ),
	.B(n1127),
	.OUT(n1804));
   XOR2 U1428 (.A(\mult_20_3/ab[5][0] ),
	.B(n1124),
	.OUT(n449));
   XOR2 U1429 (.A(\mult_20_3/ab[4][0] ),
	.B(n1122),
	.OUT(n1806));
   XOR2 U1430 (.A(\mult_20_3/ab[3][0] ),
	.B(n1118),
	.OUT(n450));
   XOR2 U1431 (.A(n1119),
	.B(\mult_20_3/ab[2][0] ),
	.OUT(n1807));
   XOR2 U1432 (.A(n1153),
	.B(n1154),
	.OUT(n1981));
   XOR2 U1433 (.A(n1160),
	.B(n1161),
	.OUT(n1982));
   XOR2 U1434 (.A(n1177),
	.B(n1983),
	.OUT(n468));
   XOR2 U1435 (.A(n1984),
	.B(\mult_20_2/ab[2][6] ),
	.OUT(n452));
   XOR2 U1436 (.A(n1185),
	.B(n1170),
	.OUT(n1985));
   XOR2 U1437 (.A(\mult_20_2/ab[4][4] ),
	.B(n1174),
	.OUT(n459));
   XOR2 U1438 (.A(\mult_20_2/ab[5][3] ),
	.B(n1176),
	.OUT(n1986));
   XOR2 U1439 (.A(\mult_20_2/ab[4][5] ),
	.B(n1183),
	.OUT(n471));
   XOR2 U1440 (.A(\mult_20_2/ab[5][4] ),
	.B(n1188),
	.OUT(n1987));
   XOR2 U1441 (.A(\mult_20_2/ab[6][3] ),
	.B(n1191),
	.OUT(n474));
   XOR2 U1442 (.A(n1988),
	.B(n1237),
	.OUT(n477));
   XOR2 U1443 (.A(\mult_20_2/ab[6][4] ),
	.B(n1197),
	.OUT(n1989));
   XOR2 U1444 (.A(\mult_20_2/ab[7][3] ),
	.B(n1199),
	.OUT(n479));
   XOR2 U1445 (.A(\mult_20_2/ab[3][2] ),
	.B(n1145),
	.OUT(n1990));
   XOR2 U1446 (.A(\mult_20_2/ab[4][2] ),
	.B(n1150),
	.OUT(n485));
   XOR2 U1447 (.A(\mult_20_2/ab[5][2] ),
	.B(n1157),
	.OUT(n1991));
   XOR2 U1448 (.A(\mult_20_2/ab[6][2] ),
	.B(n1167),
	.OUT(n488));
   XOR2 U1449 (.A(\mult_20_2/ab[7][2] ),
	.B(n1179),
	.OUT(n1992));
   XOR2 U1450 (.A(n1206),
	.B(n1203),
	.OUT(n1993));
   XOR2 U1451 (.A(\mult_20_2/ab[4][1] ),
	.B(n1207),
	.OUT(n494));
   XOR2 U1452 (.A(\mult_20_2/ab[5][1] ),
	.B(n1209),
	.OUT(n1994));
   XOR2 U1453 (.A(\mult_20_2/ab[6][1] ),
	.B(n1212),
	.OUT(n497));
   XOR2 U1454 (.A(\mult_20_2/ab[7][1] ),
	.B(n1215),
	.OUT(n1995));
   XOR2 U1455 (.A(\mult_20_2/ab[6][5] ),
	.B(n1236),
	.OUT(n500));
   XOR2 U1456 (.A(\mult_20_2/ab[7][5] ),
	.B(n1240),
	.OUT(n502));
   XOR2 U1457 (.A(\mult_20_2/ab[7][4] ),
	.B(n1242),
	.OUT(n1996));
   XOR2 U1458 (.A(\mult_20_2/ab[7][0] ),
	.B(n1229),
	.OUT(n503));
   XOR2 U1459 (.A(\mult_20_2/ab[6][0] ),
	.B(n1227),
	.OUT(n1809));
   XOR2 U1460 (.A(\mult_20_2/ab[5][0] ),
	.B(n1224),
	.OUT(n504));
   XOR2 U1461 (.A(\mult_20_2/ab[4][0] ),
	.B(n1222),
	.OUT(n1811));
   XOR2 U1462 (.A(\mult_20_2/ab[3][0] ),
	.B(n1218),
	.OUT(n505));
   XOR2 U1463 (.A(n1219),
	.B(\mult_20_2/ab[2][0] ),
	.OUT(n1812));
   XOR2 U1464 (.A(n1253),
	.B(n1254),
	.OUT(n1997));
   XOR2 U1465 (.A(n1260),
	.B(n1261),
	.OUT(n1998));
   XOR2 U1466 (.A(n1277),
	.B(n1999),
	.OUT(n523));
   XOR2 U1467 (.A(n2000),
	.B(\mult_20/ab[2][6] ),
	.OUT(n507));
   XOR2 U1468 (.A(n1285),
	.B(n1270),
	.OUT(n2001));
   XOR2 U1469 (.A(\mult_20/ab[4][4] ),
	.B(n1274),
	.OUT(n514));
   XOR2 U1470 (.A(\mult_20/ab[5][3] ),
	.B(n1276),
	.OUT(n2002));
   XOR2 U1471 (.A(\mult_20/ab[4][5] ),
	.B(n1283),
	.OUT(n526));
   XOR2 U1472 (.A(\mult_20/ab[5][4] ),
	.B(n1288),
	.OUT(n2003));
   XOR2 U1473 (.A(\mult_20/ab[6][3] ),
	.B(n1291),
	.OUT(n529));
   XOR2 U1474 (.A(n2004),
	.B(n1337),
	.OUT(n532));
   XOR2 U1475 (.A(\mult_20/ab[6][4] ),
	.B(n1297),
	.OUT(n2005));
   XOR2 U1476 (.A(\mult_20/ab[7][3] ),
	.B(n1299),
	.OUT(n534));
   XOR2 U1477 (.A(\mult_20/ab[3][2] ),
	.B(n1245),
	.OUT(n2006));
   XOR2 U1478 (.A(\mult_20/ab[4][2] ),
	.B(n1250),
	.OUT(n540));
   XOR2 U1479 (.A(\mult_20/ab[5][2] ),
	.B(n1257),
	.OUT(n2007));
   XOR2 U1480 (.A(\mult_20/ab[6][2] ),
	.B(n1267),
	.OUT(n543));
   XOR2 U1481 (.A(\mult_20/ab[7][2] ),
	.B(n1279),
	.OUT(n2008));
   XOR2 U1482 (.A(n1306),
	.B(n1303),
	.OUT(n2009));
   XOR2 U1483 (.A(\mult_20/ab[4][1] ),
	.B(n1307),
	.OUT(n549));
   XOR2 U1484 (.A(\mult_20/ab[5][1] ),
	.B(n1309),
	.OUT(n2010));
   XOR2 U1485 (.A(\mult_20/ab[6][1] ),
	.B(n1312),
	.OUT(n552));
   XOR2 U1486 (.A(\mult_20/ab[7][1] ),
	.B(n1315),
	.OUT(n2011));
   XOR2 U1487 (.A(\mult_20/ab[6][5] ),
	.B(n1336),
	.OUT(n555));
   XOR2 U1488 (.A(\mult_20/ab[7][5] ),
	.B(n1340),
	.OUT(n557));
   XOR2 U1489 (.A(\mult_20/ab[7][4] ),
	.B(n1342),
	.OUT(n2012));
   XOR2 U1490 (.A(\mult_20/ab[7][0] ),
	.B(n1329),
	.OUT(n558));
   XOR2 U1491 (.A(\mult_20/ab[6][0] ),
	.B(n1327),
	.OUT(n1814));
   XOR2 U1492 (.A(\mult_20/ab[5][0] ),
	.B(n1324),
	.OUT(n559));
   XOR2 U1493 (.A(\mult_20/ab[4][0] ),
	.B(n1322),
	.OUT(n1816));
   XOR2 U1494 (.A(\mult_20/ab[3][0] ),
	.B(n1318),
	.OUT(n560));
   XOR2 U1495 (.A(n1319),
	.B(\mult_20/ab[2][0] ),
	.OUT(n1817));
   XOR2 U1496 (.A(n1353),
	.B(n1354),
	.OUT(n2013));
   XOR2 U1497 (.A(n1360),
	.B(n1361),
	.OUT(n2014));
   XOR2 U1498 (.A(n1377),
	.B(n2015),
	.OUT(n578));
   XOR2 U1499 (.A(n2016),
	.B(\mult_19_3/ab[2][6] ),
	.OUT(n562));
   XOR2 U1500 (.A(n1385),
	.B(n1370),
	.OUT(n2017));
   XOR2 U1501 (.A(\mult_19_3/ab[4][4] ),
	.B(n1374),
	.OUT(n569));
   XOR2 U1502 (.A(\mult_19_3/ab[5][3] ),
	.B(n1376),
	.OUT(n2018));
   XOR2 U1503 (.A(\mult_19_3/ab[4][5] ),
	.B(n1383),
	.OUT(n581));
   XOR2 U1504 (.A(\mult_19_3/ab[5][4] ),
	.B(n1388),
	.OUT(n2019));
   XOR2 U1505 (.A(\mult_19_3/ab[6][3] ),
	.B(n1391),
	.OUT(n584));
   XOR2 U1506 (.A(n2020),
	.B(n1437),
	.OUT(n587));
   XOR2 U1507 (.A(\mult_19_3/ab[6][4] ),
	.B(n1397),
	.OUT(n2021));
   XOR2 U1508 (.A(\mult_19_3/ab[7][3] ),
	.B(n1399),
	.OUT(n589));
   XOR2 U1509 (.A(\mult_19_3/ab[3][2] ),
	.B(n1345),
	.OUT(n2022));
   XOR2 U1510 (.A(\mult_19_3/ab[4][2] ),
	.B(n1350),
	.OUT(n595));
   XOR2 U1511 (.A(\mult_19_3/ab[5][2] ),
	.B(n1357),
	.OUT(n2023));
   XOR2 U1512 (.A(\mult_19_3/ab[6][2] ),
	.B(n1367),
	.OUT(n598));
   XOR2 U1513 (.A(\mult_19_3/ab[7][2] ),
	.B(n1379),
	.OUT(n2024));
   XOR2 U1514 (.A(n1406),
	.B(n1403),
	.OUT(n2025));
   XOR2 U1515 (.A(\mult_19_3/ab[4][1] ),
	.B(n1407),
	.OUT(n604));
   XOR2 U1516 (.A(\mult_19_3/ab[5][1] ),
	.B(n1409),
	.OUT(n2026));
   XOR2 U1517 (.A(\mult_19_3/ab[6][1] ),
	.B(n1412),
	.OUT(n607));
   XOR2 U1518 (.A(\mult_19_3/ab[7][1] ),
	.B(n1415),
	.OUT(n2027));
   XOR2 U1519 (.A(\mult_19_3/ab[6][5] ),
	.B(n1436),
	.OUT(n610));
   XOR2 U1520 (.A(\mult_19_3/ab[7][5] ),
	.B(n1440),
	.OUT(n612));
   XOR2 U1521 (.A(\mult_19_3/ab[7][4] ),
	.B(n1442),
	.OUT(n2028));
   XOR2 U1522 (.A(\mult_19_3/ab[7][0] ),
	.B(n1429),
	.OUT(n613));
   XOR2 U1523 (.A(\mult_19_3/ab[6][0] ),
	.B(n1427),
	.OUT(n1819));
   XOR2 U1524 (.A(\mult_19_3/ab[5][0] ),
	.B(n1424),
	.OUT(n614));
   XOR2 U1525 (.A(\mult_19_3/ab[4][0] ),
	.B(n1422),
	.OUT(n1821));
   XOR2 U1526 (.A(\mult_19_3/ab[3][0] ),
	.B(n1418),
	.OUT(n615));
   XOR2 U1527 (.A(n1419),
	.B(\mult_19_3/ab[2][0] ),
	.OUT(n1822));
   XOR2 U1528 (.A(n1453),
	.B(n1454),
	.OUT(n2029));
   XOR2 U1529 (.A(n1460),
	.B(n1461),
	.OUT(n2030));
   XOR2 U1530 (.A(n1477),
	.B(n2031),
	.OUT(n633));
   XOR2 U1531 (.A(n2032),
	.B(\mult_19_2/ab[2][6] ),
	.OUT(n617));
   XOR2 U1532 (.A(n1485),
	.B(n1470),
	.OUT(n2033));
   XOR2 U1533 (.A(\mult_19_2/ab[4][4] ),
	.B(n1474),
	.OUT(n624));
   XOR2 U1534 (.A(\mult_19_2/ab[5][3] ),
	.B(n1476),
	.OUT(n2034));
   XOR2 U1535 (.A(\mult_19_2/ab[4][5] ),
	.B(n1483),
	.OUT(n636));
   XOR2 U1536 (.A(\mult_19_2/ab[5][4] ),
	.B(n1488),
	.OUT(n2035));
   XOR2 U1537 (.A(\mult_19_2/ab[6][3] ),
	.B(n1491),
	.OUT(n639));
   XOR2 U1538 (.A(n2036),
	.B(n1537),
	.OUT(n642));
   XOR2 U1539 (.A(\mult_19_2/ab[6][4] ),
	.B(n1497),
	.OUT(n2037));
   XOR2 U1540 (.A(\mult_19_2/ab[7][3] ),
	.B(n1499),
	.OUT(n644));
   XOR2 U1541 (.A(\mult_19_2/ab[3][2] ),
	.B(n1445),
	.OUT(n2038));
   XOR2 U1542 (.A(\mult_19_2/ab[4][2] ),
	.B(n1450),
	.OUT(n650));
   XOR2 U1543 (.A(\mult_19_2/ab[5][2] ),
	.B(n1457),
	.OUT(n2039));
   XOR2 U1544 (.A(\mult_19_2/ab[6][2] ),
	.B(n1467),
	.OUT(n653));
   XOR2 U1545 (.A(\mult_19_2/ab[7][2] ),
	.B(n1479),
	.OUT(n2040));
   XOR2 U1546 (.A(n1506),
	.B(n1503),
	.OUT(n2041));
   XOR2 U1547 (.A(\mult_19_2/ab[4][1] ),
	.B(n1507),
	.OUT(n659));
   XOR2 U1548 (.A(\mult_19_2/ab[5][1] ),
	.B(n1509),
	.OUT(n2042));
   XOR2 U1549 (.A(\mult_19_2/ab[6][1] ),
	.B(n1512),
	.OUT(n662));
   XOR2 U1550 (.A(\mult_19_2/ab[7][1] ),
	.B(n1515),
	.OUT(n2043));
   XOR2 U1551 (.A(\mult_19_2/ab[6][5] ),
	.B(n1536),
	.OUT(n665));
   XOR2 U1552 (.A(\mult_19_2/ab[7][5] ),
	.B(n1540),
	.OUT(n667));
   XOR2 U1553 (.A(\mult_19_2/ab[7][4] ),
	.B(n1542),
	.OUT(n2044));
   XOR2 U1554 (.A(\mult_19_2/ab[7][0] ),
	.B(n1529),
	.OUT(n668));
   XOR2 U1555 (.A(\mult_19_2/ab[6][0] ),
	.B(n1527),
	.OUT(n1824));
   XOR2 U1556 (.A(\mult_19_2/ab[5][0] ),
	.B(n1524),
	.OUT(n669));
   XOR2 U1557 (.A(\mult_19_2/ab[4][0] ),
	.B(n1522),
	.OUT(n1826));
   XOR2 U1558 (.A(\mult_19_2/ab[3][0] ),
	.B(n1518),
	.OUT(n670));
   XOR2 U1559 (.A(n1519),
	.B(\mult_19_2/ab[2][0] ),
	.OUT(n1827));
   XOR2 U1560 (.A(n1553),
	.B(n1554),
	.OUT(n2045));
   XOR2 U1561 (.A(n1560),
	.B(n1561),
	.OUT(n2046));
   XOR2 U1562 (.A(n1577),
	.B(n2047),
	.OUT(n688));
   XOR2 U1563 (.A(n2048),
	.B(\mult_19/ab[2][6] ),
	.OUT(n672));
   XOR2 U1564 (.A(n1585),
	.B(n1570),
	.OUT(n2049));
   XOR2 U1565 (.A(\mult_19/ab[4][4] ),
	.B(n1574),
	.OUT(n679));
   XOR2 U1566 (.A(\mult_19/ab[5][3] ),
	.B(n1576),
	.OUT(n2050));
   XOR2 U1567 (.A(\mult_19/ab[4][5] ),
	.B(n1583),
	.OUT(n691));
   XOR2 U1568 (.A(\mult_19/ab[5][4] ),
	.B(n1588),
	.OUT(n2051));
   XOR2 U1569 (.A(\mult_19/ab[6][3] ),
	.B(n1591),
	.OUT(n694));
   XOR2 U1570 (.A(n2052),
	.B(n1637),
	.OUT(n697));
   XOR2 U1571 (.A(\mult_19/ab[6][4] ),
	.B(n1597),
	.OUT(n2053));
   XOR2 U1572 (.A(\mult_19/ab[7][3] ),
	.B(n1599),
	.OUT(n699));
   XOR2 U1573 (.A(\mult_19/ab[3][2] ),
	.B(n1545),
	.OUT(n2054));
   XOR2 U1574 (.A(\mult_19/ab[4][2] ),
	.B(n1550),
	.OUT(n705));
   XOR2 U1575 (.A(\mult_19/ab[5][2] ),
	.B(n1557),
	.OUT(n2055));
   XOR2 U1576 (.A(\mult_19/ab[6][2] ),
	.B(n1567),
	.OUT(n708));
   XOR2 U1577 (.A(\mult_19/ab[7][2] ),
	.B(n1579),
	.OUT(n2056));
   XOR2 U1578 (.A(n1606),
	.B(n1603),
	.OUT(n2057));
   XOR2 U1579 (.A(\mult_19/ab[4][1] ),
	.B(n1607),
	.OUT(n714));
   XOR2 U1580 (.A(\mult_19/ab[5][1] ),
	.B(n1609),
	.OUT(n2058));
   XOR2 U1581 (.A(\mult_19/ab[6][1] ),
	.B(n1612),
	.OUT(n717));
   XOR2 U1582 (.A(\mult_19/ab[7][1] ),
	.B(n1615),
	.OUT(n2059));
   XOR2 U1583 (.A(\mult_19/ab[6][5] ),
	.B(n1636),
	.OUT(n720));
   XOR2 U1584 (.A(\mult_19/ab[7][5] ),
	.B(n1640),
	.OUT(n722));
   XOR2 U1585 (.A(\mult_19/ab[7][4] ),
	.B(n1642),
	.OUT(n2060));
   XOR2 U1586 (.A(\mult_19/ab[7][0] ),
	.B(n1629),
	.OUT(n723));
   XOR2 U1587 (.A(\mult_19/ab[6][0] ),
	.B(n1627),
	.OUT(n1829));
   XOR2 U1588 (.A(\mult_19/ab[5][0] ),
	.B(n1624),
	.OUT(n724));
   XOR2 U1589 (.A(\mult_19/ab[4][0] ),
	.B(n1622),
	.OUT(n1831));
   XOR2 U1590 (.A(\mult_19/ab[3][0] ),
	.B(n1618),
	.OUT(n725));
   XOR2 U1591 (.A(n1619),
	.B(\mult_19/ab[2][0] ),
	.OUT(n1832));
   XOR2 U1592 (.A(N3),
	.B(N19),
	.OUT(n2061));
   XOR2 U1593 (.A(N4),
	.B(N20),
	.OUT(n2062));
   XOR2 U1594 (.A(N5),
	.B(N21),
	.OUT(n2063));
   XOR2 U1595 (.A(N6),
	.B(N22),
	.OUT(n2064));
   XOR2 U1596 (.A(N7),
	.B(N23),
	.OUT(n2065));
   XOR2 U1597 (.A(N8),
	.B(N24),
	.OUT(n2066));
   XOR2 U1598 (.A(N9),
	.B(N25),
	.OUT(n2067));
   XOR2 U1599 (.A(N10),
	.B(N26),
	.OUT(n2068));
   XOR2 U1600 (.A(N11),
	.B(N27),
	.OUT(n2069));
   XOR2 U1601 (.A(N12),
	.B(N28),
	.OUT(n2070));
   XOR2 U1602 (.A(N13),
	.B(N29),
	.OUT(n2071));
   XOR2 U1603 (.A(N14),
	.B(N30),
	.OUT(n2072));
   XOR2 U1604 (.A(N16),
	.B(N32),
	.OUT(n2073));
   XOR2 U1605 (.A(N64),
	.B(n2073),
	.OUT(n1833));
   XOR2 U1606 (.A(n203),
	.B(n209),
	.OUT(n1834));
   XOR2 U1607 (.A(n207),
	.B(n210),
	.OUT(n1835));
   XOR2 U1608 (.A(n1689),
	.B(n1690),
	.OUT(n1837));
   XOR2 U1609 (.A(N61),
	.B(n1682),
	.OUT(n1839));
   XOR2 U1610 (.A(N60),
	.B(n1678),
	.OUT(n1841));
   XOR2 U1611 (.A(N59),
	.B(n1674),
	.OUT(n1843));
   XOR2 U1612 (.A(N58),
	.B(n1670),
	.OUT(n1845));
   XOR2 U1613 (.A(N57),
	.B(n1666),
	.OUT(n1847));
   XOR2 U1614 (.A(N56),
	.B(n1662),
	.OUT(n1849));
   XOR2 U1615 (.A(n1661),
	.B(n1663),
	.OUT(n1851));
   XOR2 U1616 (.A(N54),
	.B(n1655),
	.OUT(n1853));
   XOR2 U1617 (.A(n1654),
	.B(n1652),
	.OUT(n1855));
   XOR2 U1618 (.A(N52),
	.B(n1649),
	.OUT(n1857));
   XOR2 U1619 (.A(N51),
	.B(n1646),
	.OUT(n1859));
   XOR2 U1620 (.A(n2074),
	.B(n729),
	.OUT(n1860));
   XOR2 U1621 (.A(N163),
	.B(N179),
	.OUT(n2075));
   XOR2 U1622 (.A(N164),
	.B(N180),
	.OUT(n2076));
   XOR2 U1623 (.A(N165),
	.B(N181),
	.OUT(n2077));
   XOR2 U1624 (.A(N166),
	.B(N182),
	.OUT(n2078));
   XOR2 U1625 (.A(N167),
	.B(N183),
	.OUT(n2079));
   XOR2 U1626 (.A(N168),
	.B(N184),
	.OUT(n2080));
   XOR2 U1627 (.A(N169),
	.B(N185),
	.OUT(n2081));
   XOR2 U1628 (.A(N170),
	.B(N186),
	.OUT(n2082));
   XOR2 U1629 (.A(N171),
	.B(N187),
	.OUT(n2083));
   XOR2 U1630 (.A(N172),
	.B(N188),
	.OUT(n2084));
   XOR2 U1631 (.A(N173),
	.B(N189),
	.OUT(n2085));
   XOR2 U1632 (.A(N174),
	.B(N190),
	.OUT(n2086));
   XOR2 U1633 (.A(N176),
	.B(N192),
	.OUT(n2087));
   XOR2 U1634 (.A(N224),
	.B(n2087),
	.OUT(n1861));
   XOR2 U1635 (.A(n213),
	.B(n219),
	.OUT(n1862));
   XOR2 U1636 (.A(n217),
	.B(n220),
	.OUT(n1863));
   XOR2 U1637 (.A(n1737),
	.B(n1738),
	.OUT(n1865));
   XOR2 U1638 (.A(N221),
	.B(n1730),
	.OUT(n1867));
   XOR2 U1639 (.A(N220),
	.B(n1726),
	.OUT(n1869));
   XOR2 U1640 (.A(N219),
	.B(n1722),
	.OUT(n1871));
   XOR2 U1641 (.A(N218),
	.B(n1718),
	.OUT(n1873));
   XOR2 U1642 (.A(N217),
	.B(n1714),
	.OUT(n1875));
   XOR2 U1643 (.A(N216),
	.B(n1710),
	.OUT(n1877));
   XOR2 U1644 (.A(n1709),
	.B(n1711),
	.OUT(n1879));
   XOR2 U1645 (.A(N214),
	.B(n1703),
	.OUT(n1881));
   XOR2 U1646 (.A(n1702),
	.B(n1700),
	.OUT(n1883));
   XOR2 U1647 (.A(N212),
	.B(n1697),
	.OUT(n1885));
   XOR2 U1648 (.A(N211),
	.B(n1694),
	.OUT(n1887));
   XOR2 U1649 (.A(n2088),
	.B(n735),
	.OUT(n1888));
   XOR2 U1650 (.A(N83),
	.B(N99),
	.OUT(n2089));
   XOR2 U1651 (.A(N84),
	.B(N100),
	.OUT(n2090));
   XOR2 U1652 (.A(N85),
	.B(N101),
	.OUT(n2091));
   XOR2 U1653 (.A(N86),
	.B(N102),
	.OUT(n2092));
   XOR2 U1654 (.A(N87),
	.B(N103),
	.OUT(n2093));
   XOR2 U1655 (.A(N88),
	.B(N104),
	.OUT(n2094));
   XOR2 U1656 (.A(N89),
	.B(N105),
	.OUT(n2095));
   XOR2 U1657 (.A(N90),
	.B(N106),
	.OUT(n2096));
   XOR2 U1658 (.A(N91),
	.B(N107),
	.OUT(n2097));
   XOR2 U1659 (.A(N92),
	.B(N108),
	.OUT(n2098));
   XOR2 U1660 (.A(N93),
	.B(N109),
	.OUT(n2099));
   XOR2 U1661 (.A(N94),
	.B(N110),
	.OUT(n2100));
   XOR2 U1662 (.A(N96),
	.B(N112),
	.OUT(n2101));
   XOR2 U1663 (.A(N144),
	.B(n2101),
	.OUT(n1889));
   XOR2 U1664 (.A(n223),
	.B(n229),
	.OUT(n1890));
   XOR2 U1665 (.A(n227),
	.B(n230),
	.OUT(n1891));
   XOR2 U1666 (.A(n1785),
	.B(n1786),
	.OUT(n1893));
   XOR2 U1667 (.A(N141),
	.B(n1778),
	.OUT(n1895));
   XOR2 U1668 (.A(N140),
	.B(n1774),
	.OUT(n1897));
   XOR2 U1669 (.A(N139),
	.B(n1770),
	.OUT(n1899));
   XOR2 U1670 (.A(N138),
	.B(n1766),
	.OUT(n1901));
   XOR2 U1671 (.A(N137),
	.B(n1762),
	.OUT(n1903));
   XOR2 U1672 (.A(N136),
	.B(n1758),
	.OUT(n1905));
   XOR2 U1673 (.A(n1757),
	.B(n1759),
	.OUT(n1907));
   XOR2 U1674 (.A(N134),
	.B(n1751),
	.OUT(n1909));
   XOR2 U1675 (.A(n1750),
	.B(n1748),
	.OUT(n1911));
   XOR2 U1676 (.A(N132),
	.B(n1745),
	.OUT(n1913));
   XOR2 U1677 (.A(N131),
	.B(n1742),
	.OUT(n1915));
   XOR2 U1678 (.A(n2102),
	.B(n741),
	.OUT(n1916));
   inverter U1679 (.IN(n1569),
	.OUT(n2048));
   inverter U1680 (.IN(n1559),
	.OUT(n2103));
   inverter U1681 (.IN(n1552),
	.OUT(n2104));
   inverter U1682 (.IN(n1548),
	.OUT(n2105));
   inverter U1683 (.IN(n1544),
	.OUT(n1546));
   inverter U1684 (.IN(n1602),
	.OUT(n2106));
   inverter U1685 (.IN(n1617),
	.OUT(n1619));
   inverter U1686 (.IN(n1469),
	.OUT(n2032));
   inverter U1687 (.IN(n1459),
	.OUT(n2107));
   inverter U1688 (.IN(n1452),
	.OUT(n2108));
   inverter U1689 (.IN(n1448),
	.OUT(n2109));
   inverter U1690 (.IN(n1444),
	.OUT(n1446));
   inverter U1691 (.IN(n1502),
	.OUT(n2110));
   inverter U1692 (.IN(n1517),
	.OUT(n1519));
   inverter U1693 (.IN(n1644),
	.OUT(n2111));
   inverter U1694 (.IN(n1369),
	.OUT(n2016));
   inverter U1695 (.IN(n1359),
	.OUT(n2112));
   inverter U1696 (.IN(n1352),
	.OUT(n2113));
   inverter U1697 (.IN(n1348),
	.OUT(n2114));
   inverter U1698 (.IN(n1344),
	.OUT(n1346));
   inverter U1699 (.IN(n1402),
	.OUT(n2115));
   inverter U1700 (.IN(n1417),
	.OUT(n1419));
   inverter U1701 (.IN(n1645),
	.OUT(n2074));
   inverter U1702 (.IN(n1269),
	.OUT(n2000));
   inverter U1703 (.IN(n1259),
	.OUT(n2116));
   inverter U1704 (.IN(n1252),
	.OUT(n2117));
   inverter U1705 (.IN(n1248),
	.OUT(n2118));
   inverter U1706 (.IN(n1244),
	.OUT(n1246));
   inverter U1707 (.IN(n1302),
	.OUT(n2119));
   inverter U1708 (.IN(n1317),
	.OUT(n1319));
   inverter U1709 (.IN(n1169),
	.OUT(n1984));
   inverter U1710 (.IN(n1159),
	.OUT(n2120));
   inverter U1711 (.IN(n1152),
	.OUT(n2121));
   inverter U1712 (.IN(n1148),
	.OUT(n2122));
   inverter U1713 (.IN(n1144),
	.OUT(n1146));
   inverter U1714 (.IN(n1202),
	.OUT(n2123));
   inverter U1715 (.IN(n1217),
	.OUT(n1219));
   inverter U1716 (.IN(n1740),
	.OUT(n2124));
   inverter U1717 (.IN(n1069),
	.OUT(n1968));
   inverter U1718 (.IN(n1059),
	.OUT(n2125));
   inverter U1719 (.IN(n1052),
	.OUT(n2126));
   inverter U1720 (.IN(n1048),
	.OUT(n2127));
   inverter U1721 (.IN(n1044),
	.OUT(n1046));
   inverter U1722 (.IN(n1102),
	.OUT(n2128));
   inverter U1723 (.IN(n1117),
	.OUT(n1119));
   inverter U1724 (.IN(n1741),
	.OUT(n2102));
   inverter U1725 (.IN(n969),
	.OUT(n1952));
   inverter U1726 (.IN(n959),
	.OUT(n2129));
   inverter U1727 (.IN(n952),
	.OUT(n2130));
   inverter U1728 (.IN(n948),
	.OUT(n2131));
   inverter U1729 (.IN(n944),
	.OUT(n946));
   inverter U1730 (.IN(n1002),
	.OUT(n2132));
   inverter U1731 (.IN(n1017),
	.OUT(n1019));
   inverter U1732 (.IN(n869),
	.OUT(n1936));
   inverter U1733 (.IN(n859),
	.OUT(n2133));
   inverter U1734 (.IN(n852),
	.OUT(n2134));
   inverter U1735 (.IN(n848),
	.OUT(n2135));
   inverter U1736 (.IN(n844),
	.OUT(n846));
   inverter U1737 (.IN(n902),
	.OUT(n2136));
   inverter U1738 (.IN(n917),
	.OUT(n919));
   inverter U1739 (.IN(n1692),
	.OUT(n2137));
   inverter U1740 (.IN(n769),
	.OUT(n1920));
   inverter U1741 (.IN(n759),
	.OUT(n2138));
   inverter U1742 (.IN(n752),
	.OUT(n2139));
   inverter U1743 (.IN(n748),
	.OUT(n2140));
   inverter U1744 (.IN(n744),
	.OUT(n746));
   inverter U1745 (.IN(n802),
	.OUT(n2141));
   inverter U1746 (.IN(n817),
	.OUT(n819));
   inverter U1747 (.IN(n1693),
	.OUT(n2088));
   OAI21 U1748 (.OUT(n2142),
	.C(n1920),
	.B(\mult_21_3/ab[2][6] ),
	.A(\mult_21_3/ab[1][7] ));
   AOI21 U1749 (.OUT(n2143),
	.C(n2144),
	.B(\mult_21_3/ab[1][7] ),
	.A(\mult_21_3/ab[2][6] ));
   AOI21 U1750 (.OUT(n2145),
	.C(n2143),
	.B(n781),
	.A(n782));
   AOI21 U1751 (.OUT(n2146),
	.C(n2145),
	.B(\mult_21_3/ab[2][7] ),
	.A(\mult_21_3/ab[3][6] ));
   OAI21 U1752 (.OUT(n772),
	.C(n233),
	.B(n2138),
	.A(\mult_21_3/ab[2][5] ));
   inverter U1753 (.IN(n770),
	.OUT(n784));
   OAI21 U1754 (.OUT(n786),
	.C(n231),
	.B(n770),
	.A(\mult_21_3/ab[3][5] ));
   OAI21 U1755 (.OUT(n2147),
	.C(n250),
	.B(n783),
	.A(\mult_21_3/ab[4][5] ));
   inverter U1756 (.IN(n795),
	.OUT(n837));
   OAI21 U1757 (.OUT(n763),
	.C(n234),
	.B(n2139),
	.A(\mult_21_3/ab[2][4] ));
   AOI21 U1758 (.OUT(n775),
	.C(n235),
	.B(n2148),
	.A(n760));
   AOI21 U1759 (.OUT(n790),
	.C(n238),
	.B(n774),
	.A(n773));
   OAI21 U1760 (.OUT(n798),
	.C(n249),
	.B(n2149),
	.A(\mult_21_3/ab[5][4] ));
   OAI21 U1761 (.OUT(n756),
	.C(n240),
	.B(n2140),
	.A(\mult_21_3/ab[2][3] ));
   AOI21 U1762 (.OUT(n765),
	.C(n241),
	.B(n2150),
	.A(n753));
   inverter U1763 (.IN(n764),
	.OUT(n1919));
   OAI21 U1764 (.OUT(n778),
	.C(n247),
	.B(n1919),
	.A(\mult_21_3/ab[4][3] ));
   OAI21 U1765 (.OUT(n2151),
	.C(n237),
	.B(n776),
	.A(\mult_21_3/ab[5][3] ));
   AOI21 U1766 (.OUT(n2152),
	.C(n253),
	.B(n791),
	.A(n800));
   OAI21 U1767 (.OUT(n2153),
	.C(n243),
	.B(n746),
	.A(\mult_21_3/ab[2][2] ));
   AOI21 U1768 (.OUT(n2154),
	.C(n244),
	.B(n745),
	.A(n749));
   OAI21 U1769 (.OUT(n2155),
	.C(n264),
	.B(n750),
	.A(\mult_21_3/ab[4][2] ));
   AOI21 U1770 (.OUT(n2156),
	.C(n246),
	.B(n757),
	.A(n766));
   OAI21 U1771 (.OUT(n2157),
	.C(n267),
	.B(n767),
	.A(\mult_21_3/ab[6][2] ));
   inverter U1772 (.IN(n779),
	.OUT(n2158));
   OAI21 U1773 (.OUT(n2159),
	.C(n252),
	.B(n2158),
	.A(\mult_21_3/ab[7][2] ));
   AOI21 U1774 (.OUT(n195),
	.C(n2160),
	.B(\mult_21_3/ab[7][2] ),
	.A(n2158));
   OAI21 U1775 (.OUT(n805),
	.C(n260),
	.B(n2141),
	.A(\mult_21_3/ab[2][1] ));
   AOI21 U1776 (.OUT(n808),
	.C(n261),
	.B(n2161),
	.A(n806));
   inverter U1777 (.IN(n807),
	.OUT(n2162));
   OAI21 U1778 (.OUT(n811),
	.C(n273),
	.B(n2162),
	.A(\mult_21_3/ab[4][1] ));
   OAI21 U1779 (.OUT(n2163),
	.C(n263),
	.B(n809),
	.A(\mult_21_3/ab[5][1] ));
   inverter U1780 (.IN(n812),
	.OUT(n2164));
   OAI21 U1781 (.OUT(n816),
	.C(n276),
	.B(n2164),
	.A(\mult_21_3/ab[6][1] ));
   OAI21 U1782 (.OUT(n2165),
	.C(n266),
	.B(n815),
	.A(\mult_21_3/ab[7][1] ));
   AOI21 U1783 (.OUT(n197),
	.C(n2166),
	.B(\mult_21_3/ab[7][1] ),
	.A(n815));
   OAI21 U1784 (.OUT(n2167),
	.C(n269),
	.B(n819),
	.A(\mult_21_3/ab[2][0] ));
   AOI21 U1785 (.OUT(n2168),
	.C(n270),
	.B(n818),
	.A(n821));
   OAI21 U1786 (.OUT(n2169),
	.C(n1790),
	.B(n822),
	.A(\mult_21_3/ab[4][0] ));
   AOI21 U1787 (.OUT(n2170),
	.C(n272),
	.B(n824),
	.A(n826));
   OAI21 U1788 (.OUT(n2171),
	.C(n1788),
	.B(n827),
	.A(\mult_21_3/ab[6][0] ));
   inverter U1789 (.IN(n829),
	.OUT(n2172));
   AOI21 U1790 (.OUT(n2173),
	.C(n275),
	.B(n829),
	.A(n831));
   AOI21 U1791 (.OUT(n199),
	.C(n2173),
	.B(\mult_21_3/ab[7][0] ),
	.A(n2172));
   AOI21 U1792 (.OUT(n2174),
	.C(n2146),
	.B(n793),
	.A(n794));
   AOI21 U1793 (.OUT(n2175),
	.C(n2174),
	.B(\mult_21_3/ab[3][7] ),
	.A(\mult_21_3/ab[4][6] ));
   AOI21 U1794 (.OUT(n2176),
	.C(n2175),
	.B(n833),
	.A(n832));
   AOI21 U1795 (.OUT(n2177),
	.C(n2176),
	.B(\mult_21_3/ab[5][6] ),
	.A(\mult_21_3/ab[4][7] ));
   AOI21 U1796 (.OUT(n2178),
	.C(n2177),
	.B(n835),
	.A(n834));
   AOI21 U1797 (.OUT(n2179),
	.C(n2178),
	.B(\mult_21_3/ab[6][6] ),
	.A(\mult_21_3/ab[5][7] ));
   OAI21 U1798 (.OUT(n2180),
	.C(n2181),
	.B(\mult_21_3/ab[7][6] ),
	.A(\mult_21_3/ab[6][7] ));
   AOI21 U1799 (.OUT(n186),
	.C(n2182),
	.B(\mult_21_3/ab[7][6] ),
	.A(\mult_21_3/ab[6][7] ));
   AOI21 U1800 (.OUT(n838),
	.C(n256),
	.B(n795),
	.A(n1924));
   AOI21 U1801 (.OUT(n2183),
	.C(n279),
	.B(n836),
	.A(n839));
   OAI21 U1802 (.OUT(n2184),
	.C(n281),
	.B(n840),
	.A(\mult_21_3/ab[7][5] ));
   AOI21 U1803 (.OUT(n188),
	.C(n2185),
	.B(\mult_21_3/ab[7][5] ),
	.A(n840));
   OAI21 U1804 (.OUT(n2186),
	.C(n255),
	.B(n797),
	.A(\mult_21_3/ab[6][4] ));
   inverter U1805 (.IN(n842),
	.OUT(n2187));
   OAI21 U1806 (.OUT(n2188),
	.C(n278),
	.B(n2187),
	.A(\mult_21_3/ab[7][4] ));
   OAI21 U1807 (.OUT(n191),
	.C(n2188),
	.B(n2189),
	.A(n842));
   OAI21 U1808 (.OUT(n2190),
	.C(n2191),
	.B(n799),
	.A(\mult_21_3/ab[7][3] ));
   AOI21 U1809 (.OUT(n193),
	.C(n2192),
	.B(\mult_21_3/ab[7][3] ),
	.A(n799));
   OAI21 U1810 (.OUT(n2193),
	.C(n1936),
	.B(\mult_21_2/ab[2][6] ),
	.A(\mult_21_2/ab[1][7] ));
   AOI21 U1811 (.OUT(n2194),
	.C(n2195),
	.B(\mult_21_2/ab[1][7] ),
	.A(\mult_21_2/ab[2][6] ));
   AOI21 U1812 (.OUT(n2196),
	.C(n2194),
	.B(n881),
	.A(n882));
   AOI21 U1813 (.OUT(n2197),
	.C(n2196),
	.B(\mult_21_2/ab[2][7] ),
	.A(\mult_21_2/ab[3][6] ));
   OAI21 U1814 (.OUT(n872),
	.C(n288),
	.B(n2133),
	.A(\mult_21_2/ab[2][5] ));
   inverter U1815 (.IN(n870),
	.OUT(n884));
   OAI21 U1816 (.OUT(n886),
	.C(n286),
	.B(n870),
	.A(\mult_21_2/ab[3][5] ));
   OAI21 U1817 (.OUT(n2198),
	.C(n305),
	.B(n883),
	.A(\mult_21_2/ab[4][5] ));
   inverter U1818 (.IN(n895),
	.OUT(n937));
   OAI21 U1819 (.OUT(n863),
	.C(n289),
	.B(n2134),
	.A(\mult_21_2/ab[2][4] ));
   AOI21 U1820 (.OUT(n875),
	.C(n290),
	.B(n2199),
	.A(n860));
   AOI21 U1821 (.OUT(n890),
	.C(n293),
	.B(n874),
	.A(n873));
   OAI21 U1822 (.OUT(n898),
	.C(n304),
	.B(n2200),
	.A(\mult_21_2/ab[5][4] ));
   OAI21 U1823 (.OUT(n856),
	.C(n295),
	.B(n2135),
	.A(\mult_21_2/ab[2][3] ));
   AOI21 U1824 (.OUT(n865),
	.C(n296),
	.B(n2201),
	.A(n853));
   inverter U1825 (.IN(n864),
	.OUT(n1935));
   OAI21 U1826 (.OUT(n878),
	.C(n302),
	.B(n1935),
	.A(\mult_21_2/ab[4][3] ));
   OAI21 U1827 (.OUT(n2202),
	.C(n292),
	.B(n876),
	.A(\mult_21_2/ab[5][3] ));
   AOI21 U1828 (.OUT(n2203),
	.C(n308),
	.B(n891),
	.A(n900));
   OAI21 U1829 (.OUT(n2204),
	.C(n298),
	.B(n846),
	.A(\mult_21_2/ab[2][2] ));
   AOI21 U1830 (.OUT(n2205),
	.C(n299),
	.B(n845),
	.A(n849));
   OAI21 U1831 (.OUT(n2206),
	.C(n319),
	.B(n850),
	.A(\mult_21_2/ab[4][2] ));
   AOI21 U1832 (.OUT(n2207),
	.C(n301),
	.B(n857),
	.A(n866));
   OAI21 U1833 (.OUT(n2208),
	.C(n322),
	.B(n867),
	.A(\mult_21_2/ab[6][2] ));
   inverter U1834 (.IN(n879),
	.OUT(n2209));
   OAI21 U1835 (.OUT(n2210),
	.C(n307),
	.B(n2209),
	.A(\mult_21_2/ab[7][2] ));
   AOI21 U1836 (.OUT(n180),
	.C(n2211),
	.B(\mult_21_2/ab[7][2] ),
	.A(n2209));
   OAI21 U1837 (.OUT(n905),
	.C(n315),
	.B(n2136),
	.A(\mult_21_2/ab[2][1] ));
   AOI21 U1838 (.OUT(n908),
	.C(n316),
	.B(n2212),
	.A(n906));
   inverter U1839 (.IN(n907),
	.OUT(n2213));
   OAI21 U1840 (.OUT(n911),
	.C(n328),
	.B(n2213),
	.A(\mult_21_2/ab[4][1] ));
   OAI21 U1841 (.OUT(n2214),
	.C(n318),
	.B(n909),
	.A(\mult_21_2/ab[5][1] ));
   inverter U1842 (.IN(n912),
	.OUT(n2215));
   OAI21 U1843 (.OUT(n916),
	.C(n331),
	.B(n2215),
	.A(\mult_21_2/ab[6][1] ));
   OAI21 U1844 (.OUT(n2216),
	.C(n321),
	.B(n915),
	.A(\mult_21_2/ab[7][1] ));
   AOI21 U1845 (.OUT(n182),
	.C(n2217),
	.B(\mult_21_2/ab[7][1] ),
	.A(n915));
   OAI21 U1846 (.OUT(n2218),
	.C(n324),
	.B(n919),
	.A(\mult_21_2/ab[2][0] ));
   AOI21 U1847 (.OUT(n2219),
	.C(n325),
	.B(n918),
	.A(n921));
   OAI21 U1848 (.OUT(n2220),
	.C(n1795),
	.B(n922),
	.A(\mult_21_2/ab[4][0] ));
   AOI21 U1849 (.OUT(n2221),
	.C(n327),
	.B(n924),
	.A(n926));
   OAI21 U1850 (.OUT(n2222),
	.C(n1793),
	.B(n927),
	.A(\mult_21_2/ab[6][0] ));
   inverter U1851 (.IN(n929),
	.OUT(n2223));
   AOI21 U1852 (.OUT(n2224),
	.C(n330),
	.B(n929),
	.A(n931));
   AOI21 U1853 (.OUT(n184),
	.C(n2224),
	.B(\mult_21_2/ab[7][0] ),
	.A(n2223));
   AOI21 U1854 (.OUT(n2225),
	.C(n2197),
	.B(n893),
	.A(n894));
   AOI21 U1855 (.OUT(n2226),
	.C(n2225),
	.B(\mult_21_2/ab[3][7] ),
	.A(\mult_21_2/ab[4][6] ));
   AOI21 U1856 (.OUT(n2227),
	.C(n2226),
	.B(n933),
	.A(n932));
   AOI21 U1857 (.OUT(n2228),
	.C(n2227),
	.B(\mult_21_2/ab[5][6] ),
	.A(\mult_21_2/ab[4][7] ));
   AOI21 U1858 (.OUT(n2229),
	.C(n2228),
	.B(n935),
	.A(n934));
   AOI21 U1859 (.OUT(n2230),
	.C(n2229),
	.B(\mult_21_2/ab[6][6] ),
	.A(\mult_21_2/ab[5][7] ));
   OAI21 U1860 (.OUT(n2231),
	.C(n2232),
	.B(\mult_21_2/ab[7][6] ),
	.A(\mult_21_2/ab[6][7] ));
   AOI21 U1861 (.OUT(n171),
	.C(n2233),
	.B(\mult_21_2/ab[7][6] ),
	.A(\mult_21_2/ab[6][7] ));
   AOI21 U1862 (.OUT(n938),
	.C(n311),
	.B(n895),
	.A(n1940));
   AOI21 U1863 (.OUT(n2234),
	.C(n334),
	.B(n936),
	.A(n939));
   OAI21 U1864 (.OUT(n2235),
	.C(n336),
	.B(n940),
	.A(\mult_21_2/ab[7][5] ));
   AOI21 U1865 (.OUT(n173),
	.C(n2236),
	.B(\mult_21_2/ab[7][5] ),
	.A(n940));
   OAI21 U1866 (.OUT(n2237),
	.C(n310),
	.B(n897),
	.A(\mult_21_2/ab[6][4] ));
   inverter U1867 (.IN(n942),
	.OUT(n2238));
   OAI21 U1868 (.OUT(n2239),
	.C(n333),
	.B(n2238),
	.A(\mult_21_2/ab[7][4] ));
   OAI21 U1869 (.OUT(n176),
	.C(n2239),
	.B(n2240),
	.A(n942));
   OAI21 U1870 (.OUT(n2241),
	.C(n2242),
	.B(n899),
	.A(\mult_21_2/ab[7][3] ));
   AOI21 U1871 (.OUT(n178),
	.C(n2243),
	.B(\mult_21_2/ab[7][3] ),
	.A(n899));
   OAI21 U1872 (.OUT(n2244),
	.C(n1952),
	.B(\mult_21/ab[2][6] ),
	.A(\mult_21/ab[1][7] ));
   AOI21 U1873 (.OUT(n2245),
	.C(n2246),
	.B(\mult_21/ab[1][7] ),
	.A(\mult_21/ab[2][6] ));
   AOI21 U1874 (.OUT(n2247),
	.C(n2245),
	.B(n981),
	.A(n982));
   AOI21 U1875 (.OUT(n2248),
	.C(n2247),
	.B(\mult_21/ab[2][7] ),
	.A(\mult_21/ab[3][6] ));
   OAI21 U1876 (.OUT(n972),
	.C(n343),
	.B(n2129),
	.A(\mult_21/ab[2][5] ));
   inverter U1877 (.IN(n970),
	.OUT(n984));
   OAI21 U1878 (.OUT(n986),
	.C(n341),
	.B(n970),
	.A(\mult_21/ab[3][5] ));
   OAI21 U1879 (.OUT(n2249),
	.C(n360),
	.B(n983),
	.A(\mult_21/ab[4][5] ));
   inverter U1880 (.IN(n995),
	.OUT(n1037));
   OAI21 U1881 (.OUT(n963),
	.C(n344),
	.B(n2130),
	.A(\mult_21/ab[2][4] ));
   AOI21 U1882 (.OUT(n975),
	.C(n345),
	.B(n2250),
	.A(n960));
   AOI21 U1883 (.OUT(n990),
	.C(n348),
	.B(n974),
	.A(n973));
   OAI21 U1884 (.OUT(n998),
	.C(n359),
	.B(n2251),
	.A(\mult_21/ab[5][4] ));
   OAI21 U1885 (.OUT(n956),
	.C(n350),
	.B(n2131),
	.A(\mult_21/ab[2][3] ));
   AOI21 U1886 (.OUT(n965),
	.C(n351),
	.B(n2252),
	.A(n953));
   inverter U1887 (.IN(n964),
	.OUT(n1951));
   OAI21 U1888 (.OUT(n978),
	.C(n357),
	.B(n1951),
	.A(\mult_21/ab[4][3] ));
   OAI21 U1889 (.OUT(n2253),
	.C(n347),
	.B(n976),
	.A(\mult_21/ab[5][3] ));
   AOI21 U1890 (.OUT(n2254),
	.C(n363),
	.B(n991),
	.A(n1000));
   OAI21 U1891 (.OUT(n2255),
	.C(n353),
	.B(n946),
	.A(\mult_21/ab[2][2] ));
   AOI21 U1892 (.OUT(n2256),
	.C(n354),
	.B(n945),
	.A(n949));
   OAI21 U1893 (.OUT(n2257),
	.C(n374),
	.B(n950),
	.A(\mult_21/ab[4][2] ));
   AOI21 U1894 (.OUT(n2258),
	.C(n356),
	.B(n957),
	.A(n966));
   OAI21 U1895 (.OUT(n2259),
	.C(n377),
	.B(n967),
	.A(\mult_21/ab[6][2] ));
   inverter U1896 (.IN(n979),
	.OUT(n2260));
   OAI21 U1897 (.OUT(n2261),
	.C(n362),
	.B(n2260),
	.A(\mult_21/ab[7][2] ));
   AOI21 U1898 (.OUT(n165),
	.C(n2262),
	.B(\mult_21/ab[7][2] ),
	.A(n2260));
   OAI21 U1899 (.OUT(n1005),
	.C(n370),
	.B(n2132),
	.A(\mult_21/ab[2][1] ));
   AOI21 U1900 (.OUT(n1008),
	.C(n371),
	.B(n2263),
	.A(n1006));
   inverter U1901 (.IN(n1007),
	.OUT(n2264));
   OAI21 U1902 (.OUT(n1011),
	.C(n383),
	.B(n2264),
	.A(\mult_21/ab[4][1] ));
   OAI21 U1903 (.OUT(n2265),
	.C(n373),
	.B(n1009),
	.A(\mult_21/ab[5][1] ));
   inverter U1904 (.IN(n1012),
	.OUT(n2266));
   OAI21 U1905 (.OUT(n1016),
	.C(n386),
	.B(n2266),
	.A(\mult_21/ab[6][1] ));
   OAI21 U1906 (.OUT(n2267),
	.C(n376),
	.B(n1015),
	.A(\mult_21/ab[7][1] ));
   AOI21 U1907 (.OUT(n167),
	.C(n2268),
	.B(\mult_21/ab[7][1] ),
	.A(n1015));
   OAI21 U1908 (.OUT(n2269),
	.C(n379),
	.B(n1019),
	.A(\mult_21/ab[2][0] ));
   AOI21 U1909 (.OUT(n2270),
	.C(n380),
	.B(n1018),
	.A(n1021));
   OAI21 U1910 (.OUT(n2271),
	.C(n1800),
	.B(n1022),
	.A(\mult_21/ab[4][0] ));
   AOI21 U1911 (.OUT(n2272),
	.C(n382),
	.B(n1024),
	.A(n1026));
   OAI21 U1912 (.OUT(n2273),
	.C(n1798),
	.B(n1027),
	.A(\mult_21/ab[6][0] ));
   inverter U1913 (.IN(n1029),
	.OUT(n2274));
   AOI21 U1914 (.OUT(n2275),
	.C(n385),
	.B(n1029),
	.A(n1031));
   AOI21 U1915 (.OUT(n169),
	.C(n2275),
	.B(\mult_21/ab[7][0] ),
	.A(n2274));
   AOI21 U1916 (.OUT(n2276),
	.C(n2248),
	.B(n993),
	.A(n994));
   AOI21 U1917 (.OUT(n2277),
	.C(n2276),
	.B(\mult_21/ab[3][7] ),
	.A(\mult_21/ab[4][6] ));
   AOI21 U1918 (.OUT(n2278),
	.C(n2277),
	.B(n1033),
	.A(n1032));
   AOI21 U1919 (.OUT(n2279),
	.C(n2278),
	.B(\mult_21/ab[5][6] ),
	.A(\mult_21/ab[4][7] ));
   AOI21 U1920 (.OUT(n2280),
	.C(n2279),
	.B(n1035),
	.A(n1034));
   AOI21 U1921 (.OUT(n2281),
	.C(n2280),
	.B(\mult_21/ab[6][6] ),
	.A(\mult_21/ab[5][7] ));
   OAI21 U1922 (.OUT(n2282),
	.C(n2283),
	.B(\mult_21/ab[7][6] ),
	.A(\mult_21/ab[6][7] ));
   AOI21 U1923 (.OUT(n156),
	.C(n2284),
	.B(\mult_21/ab[7][6] ),
	.A(\mult_21/ab[6][7] ));
   AOI21 U1924 (.OUT(n1038),
	.C(n366),
	.B(n995),
	.A(n1956));
   AOI21 U1925 (.OUT(n2285),
	.C(n389),
	.B(n1036),
	.A(n1039));
   OAI21 U1926 (.OUT(n2286),
	.C(n391),
	.B(n1040),
	.A(\mult_21/ab[7][5] ));
   AOI21 U1927 (.OUT(n158),
	.C(n2287),
	.B(\mult_21/ab[7][5] ),
	.A(n1040));
   OAI21 U1928 (.OUT(n2288),
	.C(n365),
	.B(n997),
	.A(\mult_21/ab[6][4] ));
   inverter U1929 (.IN(n1042),
	.OUT(n2289));
   OAI21 U1930 (.OUT(n2290),
	.C(n388),
	.B(n2289),
	.A(\mult_21/ab[7][4] ));
   OAI21 U1931 (.OUT(n161),
	.C(n2290),
	.B(n2291),
	.A(n1042));
   OAI21 U1932 (.OUT(n2292),
	.C(n2293),
	.B(n999),
	.A(\mult_21/ab[7][3] ));
   AOI21 U1933 (.OUT(n163),
	.C(n2294),
	.B(\mult_21/ab[7][3] ),
	.A(n999));
   OAI21 U1934 (.OUT(n2295),
	.C(n1968),
	.B(\mult_20_3/ab[2][6] ),
	.A(\mult_20_3/ab[1][7] ));
   AOI21 U1935 (.OUT(n2296),
	.C(n2297),
	.B(\mult_20_3/ab[1][7] ),
	.A(\mult_20_3/ab[2][6] ));
   AOI21 U1936 (.OUT(n2298),
	.C(n2296),
	.B(n1081),
	.A(n1082));
   AOI21 U1937 (.OUT(n2299),
	.C(n2298),
	.B(\mult_20_3/ab[2][7] ),
	.A(\mult_20_3/ab[3][6] ));
   OAI21 U1938 (.OUT(n1072),
	.C(n398),
	.B(n2125),
	.A(\mult_20_3/ab[2][5] ));
   inverter U1939 (.IN(n1070),
	.OUT(n1084));
   OAI21 U1940 (.OUT(n1086),
	.C(n396),
	.B(n1070),
	.A(\mult_20_3/ab[3][5] ));
   OAI21 U1941 (.OUT(n2300),
	.C(n415),
	.B(n1083),
	.A(\mult_20_3/ab[4][5] ));
   inverter U1942 (.IN(n1095),
	.OUT(n1137));
   OAI21 U1943 (.OUT(n1063),
	.C(n399),
	.B(n2126),
	.A(\mult_20_3/ab[2][4] ));
   AOI21 U1944 (.OUT(n1075),
	.C(n400),
	.B(n2301),
	.A(n1060));
   AOI21 U1945 (.OUT(n1090),
	.C(n403),
	.B(n1074),
	.A(n1073));
   OAI21 U1946 (.OUT(n1098),
	.C(n414),
	.B(n2302),
	.A(\mult_20_3/ab[5][4] ));
   OAI21 U1947 (.OUT(n1056),
	.C(n405),
	.B(n2127),
	.A(\mult_20_3/ab[2][3] ));
   AOI21 U1948 (.OUT(n1065),
	.C(n406),
	.B(n2303),
	.A(n1053));
   inverter U1949 (.IN(n1064),
	.OUT(n1967));
   OAI21 U1950 (.OUT(n1078),
	.C(n412),
	.B(n1967),
	.A(\mult_20_3/ab[4][3] ));
   OAI21 U1951 (.OUT(n2304),
	.C(n402),
	.B(n1076),
	.A(\mult_20_3/ab[5][3] ));
   AOI21 U1952 (.OUT(n2305),
	.C(n418),
	.B(n1091),
	.A(n1100));
   OAI21 U1953 (.OUT(n2306),
	.C(n408),
	.B(n1046),
	.A(\mult_20_3/ab[2][2] ));
   AOI21 U1954 (.OUT(n2307),
	.C(n409),
	.B(n1045),
	.A(n1049));
   OAI21 U1955 (.OUT(n2308),
	.C(n429),
	.B(n1050),
	.A(\mult_20_3/ab[4][2] ));
   AOI21 U1956 (.OUT(n2309),
	.C(n411),
	.B(n1057),
	.A(n1066));
   OAI21 U1957 (.OUT(n2310),
	.C(n432),
	.B(n1067),
	.A(\mult_20_3/ab[6][2] ));
   inverter U1958 (.IN(n1079),
	.OUT(n2311));
   OAI21 U1959 (.OUT(n2312),
	.C(n417),
	.B(n2311),
	.A(\mult_20_3/ab[7][2] ));
   AOI21 U1960 (.OUT(n150),
	.C(n2313),
	.B(\mult_20_3/ab[7][2] ),
	.A(n2311));
   OAI21 U1961 (.OUT(n1105),
	.C(n425),
	.B(n2128),
	.A(\mult_20_3/ab[2][1] ));
   AOI21 U1962 (.OUT(n1108),
	.C(n426),
	.B(n2314),
	.A(n1106));
   inverter U1963 (.IN(n1107),
	.OUT(n2315));
   OAI21 U1964 (.OUT(n1111),
	.C(n438),
	.B(n2315),
	.A(\mult_20_3/ab[4][1] ));
   OAI21 U1965 (.OUT(n2316),
	.C(n428),
	.B(n1109),
	.A(\mult_20_3/ab[5][1] ));
   inverter U1966 (.IN(n1112),
	.OUT(n2317));
   OAI21 U1967 (.OUT(n1116),
	.C(n441),
	.B(n2317),
	.A(\mult_20_3/ab[6][1] ));
   OAI21 U1968 (.OUT(n2318),
	.C(n431),
	.B(n1115),
	.A(\mult_20_3/ab[7][1] ));
   AOI21 U1969 (.OUT(n152),
	.C(n2319),
	.B(\mult_20_3/ab[7][1] ),
	.A(n1115));
   OAI21 U1970 (.OUT(n2320),
	.C(n434),
	.B(n1119),
	.A(\mult_20_3/ab[2][0] ));
   AOI21 U1971 (.OUT(n2321),
	.C(n435),
	.B(n1118),
	.A(n1121));
   OAI21 U1972 (.OUT(n2322),
	.C(n1805),
	.B(n1122),
	.A(\mult_20_3/ab[4][0] ));
   AOI21 U1973 (.OUT(n2323),
	.C(n437),
	.B(n1124),
	.A(n1126));
   OAI21 U1974 (.OUT(n2324),
	.C(n1803),
	.B(n1127),
	.A(\mult_20_3/ab[6][0] ));
   inverter U1975 (.IN(n1129),
	.OUT(n2325));
   AOI21 U1976 (.OUT(n2326),
	.C(n440),
	.B(n1129),
	.A(n1131));
   AOI21 U1977 (.OUT(n154),
	.C(n2326),
	.B(\mult_20_3/ab[7][0] ),
	.A(n2325));
   AOI21 U1978 (.OUT(n2327),
	.C(n2299),
	.B(n1093),
	.A(n1094));
   AOI21 U1979 (.OUT(n2328),
	.C(n2327),
	.B(\mult_20_3/ab[3][7] ),
	.A(\mult_20_3/ab[4][6] ));
   AOI21 U1980 (.OUT(n2329),
	.C(n2328),
	.B(n1133),
	.A(n1132));
   AOI21 U1981 (.OUT(n2330),
	.C(n2329),
	.B(\mult_20_3/ab[5][6] ),
	.A(\mult_20_3/ab[4][7] ));
   AOI21 U1982 (.OUT(n2331),
	.C(n2330),
	.B(n1135),
	.A(n1134));
   AOI21 U1983 (.OUT(n2332),
	.C(n2331),
	.B(\mult_20_3/ab[6][6] ),
	.A(\mult_20_3/ab[5][7] ));
   OAI21 U1984 (.OUT(n2333),
	.C(n2334),
	.B(\mult_20_3/ab[7][6] ),
	.A(\mult_20_3/ab[6][7] ));
   AOI21 U1985 (.OUT(n141),
	.C(n2335),
	.B(\mult_20_3/ab[7][6] ),
	.A(\mult_20_3/ab[6][7] ));
   AOI21 U1986 (.OUT(n1138),
	.C(n421),
	.B(n1095),
	.A(n1972));
   AOI21 U1987 (.OUT(n2336),
	.C(n444),
	.B(n1136),
	.A(n1139));
   OAI21 U1988 (.OUT(n2337),
	.C(n446),
	.B(n1140),
	.A(\mult_20_3/ab[7][5] ));
   AOI21 U1989 (.OUT(n143),
	.C(n2338),
	.B(\mult_20_3/ab[7][5] ),
	.A(n1140));
   OAI21 U1990 (.OUT(n2339),
	.C(n420),
	.B(n1097),
	.A(\mult_20_3/ab[6][4] ));
   inverter U1991 (.IN(n1142),
	.OUT(n2340));
   OAI21 U1992 (.OUT(n2341),
	.C(n443),
	.B(n2340),
	.A(\mult_20_3/ab[7][4] ));
   OAI21 U1993 (.OUT(n146),
	.C(n2341),
	.B(n2342),
	.A(n1142));
   OAI21 U1994 (.OUT(n2343),
	.C(n2344),
	.B(n1099),
	.A(\mult_20_3/ab[7][3] ));
   AOI21 U1995 (.OUT(n148),
	.C(n2345),
	.B(\mult_20_3/ab[7][3] ),
	.A(n1099));
   OAI21 U1996 (.OUT(n2346),
	.C(n1984),
	.B(\mult_20_2/ab[2][6] ),
	.A(\mult_20_2/ab[1][7] ));
   AOI21 U1997 (.OUT(n2347),
	.C(n2348),
	.B(\mult_20_2/ab[1][7] ),
	.A(\mult_20_2/ab[2][6] ));
   AOI21 U1998 (.OUT(n2349),
	.C(n2347),
	.B(n1181),
	.A(n1182));
   AOI21 U1999 (.OUT(n2350),
	.C(n2349),
	.B(\mult_20_2/ab[2][7] ),
	.A(\mult_20_2/ab[3][6] ));
   OAI21 U2000 (.OUT(n1172),
	.C(n453),
	.B(n2120),
	.A(\mult_20_2/ab[2][5] ));
   inverter U2001 (.IN(n1170),
	.OUT(n1184));
   OAI21 U2002 (.OUT(n1186),
	.C(n451),
	.B(n1170),
	.A(\mult_20_2/ab[3][5] ));
   OAI21 U2003 (.OUT(n2351),
	.C(n470),
	.B(n1183),
	.A(\mult_20_2/ab[4][5] ));
   inverter U2004 (.IN(n1195),
	.OUT(n1237));
   OAI21 U2005 (.OUT(n1163),
	.C(n454),
	.B(n2121),
	.A(\mult_20_2/ab[2][4] ));
   AOI21 U2006 (.OUT(n1175),
	.C(n455),
	.B(n2352),
	.A(n1160));
   AOI21 U2007 (.OUT(n1190),
	.C(n458),
	.B(n1174),
	.A(n1173));
   OAI21 U2008 (.OUT(n1198),
	.C(n469),
	.B(n2353),
	.A(\mult_20_2/ab[5][4] ));
   OAI21 U2009 (.OUT(n1156),
	.C(n460),
	.B(n2122),
	.A(\mult_20_2/ab[2][3] ));
   AOI21 U2010 (.OUT(n1165),
	.C(n461),
	.B(n2354),
	.A(n1153));
   inverter U2011 (.IN(n1164),
	.OUT(n1983));
   OAI21 U2012 (.OUT(n1178),
	.C(n467),
	.B(n1983),
	.A(\mult_20_2/ab[4][3] ));
   OAI21 U2013 (.OUT(n2355),
	.C(n457),
	.B(n1176),
	.A(\mult_20_2/ab[5][3] ));
   AOI21 U2014 (.OUT(n2356),
	.C(n473),
	.B(n1191),
	.A(n1200));
   OAI21 U2015 (.OUT(n2357),
	.C(n463),
	.B(n1146),
	.A(\mult_20_2/ab[2][2] ));
   AOI21 U2016 (.OUT(n2358),
	.C(n464),
	.B(n1145),
	.A(n1149));
   OAI21 U2017 (.OUT(n2359),
	.C(n484),
	.B(n1150),
	.A(\mult_20_2/ab[4][2] ));
   AOI21 U2018 (.OUT(n2360),
	.C(n466),
	.B(n1157),
	.A(n1166));
   OAI21 U2019 (.OUT(n2361),
	.C(n487),
	.B(n1167),
	.A(\mult_20_2/ab[6][2] ));
   inverter U2020 (.IN(n1179),
	.OUT(n2362));
   OAI21 U2021 (.OUT(n2363),
	.C(n472),
	.B(n2362),
	.A(\mult_20_2/ab[7][2] ));
   AOI21 U2022 (.OUT(n135),
	.C(n2364),
	.B(\mult_20_2/ab[7][2] ),
	.A(n2362));
   OAI21 U2023 (.OUT(n1205),
	.C(n480),
	.B(n2123),
	.A(\mult_20_2/ab[2][1] ));
   AOI21 U2024 (.OUT(n1208),
	.C(n481),
	.B(n2365),
	.A(n1206));
   inverter U2025 (.IN(n1207),
	.OUT(n2366));
   OAI21 U2026 (.OUT(n1211),
	.C(n493),
	.B(n2366),
	.A(\mult_20_2/ab[4][1] ));
   OAI21 U2027 (.OUT(n2367),
	.C(n483),
	.B(n1209),
	.A(\mult_20_2/ab[5][1] ));
   inverter U2028 (.IN(n1212),
	.OUT(n2368));
   OAI21 U2029 (.OUT(n1216),
	.C(n496),
	.B(n2368),
	.A(\mult_20_2/ab[6][1] ));
   OAI21 U2030 (.OUT(n2369),
	.C(n486),
	.B(n1215),
	.A(\mult_20_2/ab[7][1] ));
   AOI21 U2031 (.OUT(n137),
	.C(n2370),
	.B(\mult_20_2/ab[7][1] ),
	.A(n1215));
   OAI21 U2032 (.OUT(n2371),
	.C(n489),
	.B(n1219),
	.A(\mult_20_2/ab[2][0] ));
   AOI21 U2033 (.OUT(n2372),
	.C(n490),
	.B(n1218),
	.A(n1221));
   OAI21 U2034 (.OUT(n2373),
	.C(n1810),
	.B(n1222),
	.A(\mult_20_2/ab[4][0] ));
   AOI21 U2035 (.OUT(n2374),
	.C(n492),
	.B(n1224),
	.A(n1226));
   OAI21 U2036 (.OUT(n2375),
	.C(n1808),
	.B(n1227),
	.A(\mult_20_2/ab[6][0] ));
   inverter U2037 (.IN(n1229),
	.OUT(n2376));
   AOI21 U2038 (.OUT(n2377),
	.C(n495),
	.B(n1229),
	.A(n1231));
   AOI21 U2039 (.OUT(n139),
	.C(n2377),
	.B(\mult_20_2/ab[7][0] ),
	.A(n2376));
   AOI21 U2040 (.OUT(n2378),
	.C(n2350),
	.B(n1193),
	.A(n1194));
   AOI21 U2041 (.OUT(n2379),
	.C(n2378),
	.B(\mult_20_2/ab[3][7] ),
	.A(\mult_20_2/ab[4][6] ));
   AOI21 U2042 (.OUT(n2380),
	.C(n2379),
	.B(n1233),
	.A(n1232));
   AOI21 U2043 (.OUT(n2381),
	.C(n2380),
	.B(\mult_20_2/ab[5][6] ),
	.A(\mult_20_2/ab[4][7] ));
   AOI21 U2044 (.OUT(n2382),
	.C(n2381),
	.B(n1235),
	.A(n1234));
   AOI21 U2045 (.OUT(n2383),
	.C(n2382),
	.B(\mult_20_2/ab[6][6] ),
	.A(\mult_20_2/ab[5][7] ));
   OAI21 U2046 (.OUT(n2384),
	.C(n2385),
	.B(\mult_20_2/ab[7][6] ),
	.A(\mult_20_2/ab[6][7] ));
   AOI21 U2047 (.OUT(n126),
	.C(n2386),
	.B(\mult_20_2/ab[7][6] ),
	.A(\mult_20_2/ab[6][7] ));
   AOI21 U2048 (.OUT(n1238),
	.C(n476),
	.B(n1195),
	.A(n1988));
   AOI21 U2049 (.OUT(n2387),
	.C(n499),
	.B(n1236),
	.A(n1239));
   OAI21 U2050 (.OUT(n2388),
	.C(n501),
	.B(n1240),
	.A(\mult_20_2/ab[7][5] ));
   AOI21 U2051 (.OUT(n128),
	.C(n2389),
	.B(\mult_20_2/ab[7][5] ),
	.A(n1240));
   OAI21 U2052 (.OUT(n2390),
	.C(n475),
	.B(n1197),
	.A(\mult_20_2/ab[6][4] ));
   inverter U2053 (.IN(n1242),
	.OUT(n2391));
   OAI21 U2054 (.OUT(n2392),
	.C(n498),
	.B(n2391),
	.A(\mult_20_2/ab[7][4] ));
   OAI21 U2055 (.OUT(n131),
	.C(n2392),
	.B(n2393),
	.A(n1242));
   OAI21 U2056 (.OUT(n2394),
	.C(n2395),
	.B(n1199),
	.A(\mult_20_2/ab[7][3] ));
   AOI21 U2057 (.OUT(n133),
	.C(n2396),
	.B(\mult_20_2/ab[7][3] ),
	.A(n1199));
   OAI21 U2058 (.OUT(n2397),
	.C(n2000),
	.B(\mult_20/ab[2][6] ),
	.A(\mult_20/ab[1][7] ));
   AOI21 U2059 (.OUT(n2398),
	.C(n2399),
	.B(\mult_20/ab[1][7] ),
	.A(\mult_20/ab[2][6] ));
   AOI21 U2060 (.OUT(n2400),
	.C(n2398),
	.B(n1281),
	.A(n1282));
   AOI21 U2061 (.OUT(n2401),
	.C(n2400),
	.B(\mult_20/ab[2][7] ),
	.A(\mult_20/ab[3][6] ));
   OAI21 U2062 (.OUT(n1272),
	.C(n508),
	.B(n2116),
	.A(\mult_20/ab[2][5] ));
   inverter U2063 (.IN(n1270),
	.OUT(n1284));
   OAI21 U2064 (.OUT(n1286),
	.C(n506),
	.B(n1270),
	.A(\mult_20/ab[3][5] ));
   OAI21 U2065 (.OUT(n2402),
	.C(n525),
	.B(n1283),
	.A(\mult_20/ab[4][5] ));
   inverter U2066 (.IN(n1295),
	.OUT(n1337));
   OAI21 U2067 (.OUT(n1263),
	.C(n509),
	.B(n2117),
	.A(\mult_20/ab[2][4] ));
   AOI21 U2068 (.OUT(n1275),
	.C(n510),
	.B(n2403),
	.A(n1260));
   AOI21 U2069 (.OUT(n1290),
	.C(n513),
	.B(n1274),
	.A(n1273));
   OAI21 U2070 (.OUT(n1298),
	.C(n524),
	.B(n2404),
	.A(\mult_20/ab[5][4] ));
   OAI21 U2071 (.OUT(n1256),
	.C(n515),
	.B(n2118),
	.A(\mult_20/ab[2][3] ));
   AOI21 U2072 (.OUT(n1265),
	.C(n516),
	.B(n2405),
	.A(n1253));
   inverter U2073 (.IN(n1264),
	.OUT(n1999));
   OAI21 U2074 (.OUT(n1278),
	.C(n522),
	.B(n1999),
	.A(\mult_20/ab[4][3] ));
   OAI21 U2075 (.OUT(n2406),
	.C(n512),
	.B(n1276),
	.A(\mult_20/ab[5][3] ));
   AOI21 U2076 (.OUT(n2407),
	.C(n528),
	.B(n1291),
	.A(n1300));
   OAI21 U2077 (.OUT(n2408),
	.C(n518),
	.B(n1246),
	.A(\mult_20/ab[2][2] ));
   AOI21 U2078 (.OUT(n2409),
	.C(n519),
	.B(n1245),
	.A(n1249));
   OAI21 U2079 (.OUT(n2410),
	.C(n539),
	.B(n1250),
	.A(\mult_20/ab[4][2] ));
   AOI21 U2080 (.OUT(n2411),
	.C(n521),
	.B(n1257),
	.A(n1266));
   OAI21 U2081 (.OUT(n2412),
	.C(n542),
	.B(n1267),
	.A(\mult_20/ab[6][2] ));
   inverter U2082 (.IN(n1279),
	.OUT(n2413));
   OAI21 U2083 (.OUT(n2414),
	.C(n527),
	.B(n2413),
	.A(\mult_20/ab[7][2] ));
   AOI21 U2084 (.OUT(n120),
	.C(n2415),
	.B(\mult_20/ab[7][2] ),
	.A(n2413));
   OAI21 U2085 (.OUT(n1305),
	.C(n535),
	.B(n2119),
	.A(\mult_20/ab[2][1] ));
   AOI21 U2086 (.OUT(n1308),
	.C(n536),
	.B(n2416),
	.A(n1306));
   inverter U2087 (.IN(n1307),
	.OUT(n2417));
   OAI21 U2088 (.OUT(n1311),
	.C(n548),
	.B(n2417),
	.A(\mult_20/ab[4][1] ));
   OAI21 U2089 (.OUT(n2418),
	.C(n538),
	.B(n1309),
	.A(\mult_20/ab[5][1] ));
   inverter U2090 (.IN(n1312),
	.OUT(n2419));
   OAI21 U2091 (.OUT(n1316),
	.C(n551),
	.B(n2419),
	.A(\mult_20/ab[6][1] ));
   OAI21 U2092 (.OUT(n2420),
	.C(n541),
	.B(n1315),
	.A(\mult_20/ab[7][1] ));
   AOI21 U2093 (.OUT(n122),
	.C(n2421),
	.B(\mult_20/ab[7][1] ),
	.A(n1315));
   OAI21 U2094 (.OUT(n2422),
	.C(n544),
	.B(n1319),
	.A(\mult_20/ab[2][0] ));
   AOI21 U2095 (.OUT(n2423),
	.C(n545),
	.B(n1318),
	.A(n1321));
   OAI21 U2096 (.OUT(n2424),
	.C(n1815),
	.B(n1322),
	.A(\mult_20/ab[4][0] ));
   AOI21 U2097 (.OUT(n2425),
	.C(n547),
	.B(n1324),
	.A(n1326));
   OAI21 U2098 (.OUT(n2426),
	.C(n1813),
	.B(n1327),
	.A(\mult_20/ab[6][0] ));
   inverter U2099 (.IN(n1329),
	.OUT(n2427));
   AOI21 U2100 (.OUT(n2428),
	.C(n550),
	.B(n1329),
	.A(n1331));
   AOI21 U2101 (.OUT(n124),
	.C(n2428),
	.B(\mult_20/ab[7][0] ),
	.A(n2427));
   AOI21 U2102 (.OUT(n2429),
	.C(n2401),
	.B(n1293),
	.A(n1294));
   AOI21 U2103 (.OUT(n2430),
	.C(n2429),
	.B(\mult_20/ab[3][7] ),
	.A(\mult_20/ab[4][6] ));
   AOI21 U2104 (.OUT(n2431),
	.C(n2430),
	.B(n1333),
	.A(n1332));
   AOI21 U2105 (.OUT(n2432),
	.C(n2431),
	.B(\mult_20/ab[5][6] ),
	.A(\mult_20/ab[4][7] ));
   AOI21 U2106 (.OUT(n2433),
	.C(n2432),
	.B(n1335),
	.A(n1334));
   AOI21 U2107 (.OUT(n2434),
	.C(n2433),
	.B(\mult_20/ab[6][6] ),
	.A(\mult_20/ab[5][7] ));
   OAI21 U2108 (.OUT(n2435),
	.C(n2436),
	.B(\mult_20/ab[7][6] ),
	.A(\mult_20/ab[6][7] ));
   AOI21 U2109 (.OUT(n111),
	.C(n2437),
	.B(\mult_20/ab[7][6] ),
	.A(\mult_20/ab[6][7] ));
   AOI21 U2110 (.OUT(n1338),
	.C(n531),
	.B(n1295),
	.A(n2004));
   AOI21 U2111 (.OUT(n2438),
	.C(n554),
	.B(n1336),
	.A(n1339));
   OAI21 U2112 (.OUT(n2439),
	.C(n556),
	.B(n1340),
	.A(\mult_20/ab[7][5] ));
   AOI21 U2113 (.OUT(n113),
	.C(n2440),
	.B(\mult_20/ab[7][5] ),
	.A(n1340));
   OAI21 U2114 (.OUT(n2441),
	.C(n530),
	.B(n1297),
	.A(\mult_20/ab[6][4] ));
   inverter U2115 (.IN(n1342),
	.OUT(n2442));
   OAI21 U2116 (.OUT(n2443),
	.C(n553),
	.B(n2442),
	.A(\mult_20/ab[7][4] ));
   OAI21 U2117 (.OUT(n116),
	.C(n2443),
	.B(n2444),
	.A(n1342));
   OAI21 U2118 (.OUT(n2445),
	.C(n2446),
	.B(n1299),
	.A(\mult_20/ab[7][3] ));
   AOI21 U2119 (.OUT(n118),
	.C(n2447),
	.B(\mult_20/ab[7][3] ),
	.A(n1299));
   OAI21 U2120 (.OUT(n2448),
	.C(n2016),
	.B(\mult_19_3/ab[2][6] ),
	.A(\mult_19_3/ab[1][7] ));
   AOI21 U2121 (.OUT(n2449),
	.C(n2450),
	.B(\mult_19_3/ab[1][7] ),
	.A(\mult_19_3/ab[2][6] ));
   AOI21 U2122 (.OUT(n2451),
	.C(n2449),
	.B(n1381),
	.A(n1382));
   AOI21 U2123 (.OUT(n2452),
	.C(n2451),
	.B(\mult_19_3/ab[2][7] ),
	.A(\mult_19_3/ab[3][6] ));
   OAI21 U2124 (.OUT(n1372),
	.C(n563),
	.B(n2112),
	.A(\mult_19_3/ab[2][5] ));
   inverter U2125 (.IN(n1370),
	.OUT(n1384));
   OAI21 U2126 (.OUT(n1386),
	.C(n561),
	.B(n1370),
	.A(\mult_19_3/ab[3][5] ));
   OAI21 U2127 (.OUT(n2453),
	.C(n580),
	.B(n1383),
	.A(\mult_19_3/ab[4][5] ));
   inverter U2128 (.IN(n1395),
	.OUT(n1437));
   OAI21 U2129 (.OUT(n1363),
	.C(n564),
	.B(n2113),
	.A(\mult_19_3/ab[2][4] ));
   AOI21 U2130 (.OUT(n1375),
	.C(n565),
	.B(n2454),
	.A(n1360));
   AOI21 U2131 (.OUT(n1390),
	.C(n568),
	.B(n1374),
	.A(n1373));
   OAI21 U2132 (.OUT(n1398),
	.C(n579),
	.B(n2455),
	.A(\mult_19_3/ab[5][4] ));
   OAI21 U2133 (.OUT(n1356),
	.C(n570),
	.B(n2114),
	.A(\mult_19_3/ab[2][3] ));
   AOI21 U2134 (.OUT(n1365),
	.C(n571),
	.B(n2456),
	.A(n1353));
   inverter U2135 (.IN(n1364),
	.OUT(n2015));
   OAI21 U2136 (.OUT(n1378),
	.C(n577),
	.B(n2015),
	.A(\mult_19_3/ab[4][3] ));
   OAI21 U2137 (.OUT(n2457),
	.C(n567),
	.B(n1376),
	.A(\mult_19_3/ab[5][3] ));
   AOI21 U2138 (.OUT(n2458),
	.C(n583),
	.B(n1391),
	.A(n1400));
   OAI21 U2139 (.OUT(n2459),
	.C(n573),
	.B(n1346),
	.A(\mult_19_3/ab[2][2] ));
   AOI21 U2140 (.OUT(n2460),
	.C(n574),
	.B(n1345),
	.A(n1349));
   OAI21 U2141 (.OUT(n2461),
	.C(n594),
	.B(n1350),
	.A(\mult_19_3/ab[4][2] ));
   AOI21 U2142 (.OUT(n2462),
	.C(n576),
	.B(n1357),
	.A(n1366));
   OAI21 U2143 (.OUT(n2463),
	.C(n597),
	.B(n1367),
	.A(\mult_19_3/ab[6][2] ));
   inverter U2144 (.IN(n1379),
	.OUT(n2464));
   OAI21 U2145 (.OUT(n2465),
	.C(n582),
	.B(n2464),
	.A(\mult_19_3/ab[7][2] ));
   AOI21 U2146 (.OUT(n105),
	.C(n2466),
	.B(\mult_19_3/ab[7][2] ),
	.A(n2464));
   OAI21 U2147 (.OUT(n1405),
	.C(n590),
	.B(n2115),
	.A(\mult_19_3/ab[2][1] ));
   AOI21 U2148 (.OUT(n1408),
	.C(n591),
	.B(n2467),
	.A(n1406));
   inverter U2149 (.IN(n1407),
	.OUT(n2468));
   OAI21 U2150 (.OUT(n1411),
	.C(n603),
	.B(n2468),
	.A(\mult_19_3/ab[4][1] ));
   OAI21 U2151 (.OUT(n2469),
	.C(n593),
	.B(n1409),
	.A(\mult_19_3/ab[5][1] ));
   inverter U2152 (.IN(n1412),
	.OUT(n2470));
   OAI21 U2153 (.OUT(n1416),
	.C(n606),
	.B(n2470),
	.A(\mult_19_3/ab[6][1] ));
   OAI21 U2154 (.OUT(n2471),
	.C(n596),
	.B(n1415),
	.A(\mult_19_3/ab[7][1] ));
   AOI21 U2155 (.OUT(n107),
	.C(n2472),
	.B(\mult_19_3/ab[7][1] ),
	.A(n1415));
   OAI21 U2156 (.OUT(n2473),
	.C(n599),
	.B(n1419),
	.A(\mult_19_3/ab[2][0] ));
   AOI21 U2157 (.OUT(n2474),
	.C(n600),
	.B(n1418),
	.A(n1421));
   OAI21 U2158 (.OUT(n2475),
	.C(n1820),
	.B(n1422),
	.A(\mult_19_3/ab[4][0] ));
   AOI21 U2159 (.OUT(n2476),
	.C(n602),
	.B(n1424),
	.A(n1426));
   OAI21 U2160 (.OUT(n2477),
	.C(n1818),
	.B(n1427),
	.A(\mult_19_3/ab[6][0] ));
   inverter U2161 (.IN(n1429),
	.OUT(n2478));
   AOI21 U2162 (.OUT(n2479),
	.C(n605),
	.B(n1429),
	.A(n1431));
   AOI21 U2163 (.OUT(n109),
	.C(n2479),
	.B(\mult_19_3/ab[7][0] ),
	.A(n2478));
   AOI21 U2164 (.OUT(n2480),
	.C(n2452),
	.B(n1393),
	.A(n1394));
   AOI21 U2165 (.OUT(n2481),
	.C(n2480),
	.B(\mult_19_3/ab[3][7] ),
	.A(\mult_19_3/ab[4][6] ));
   AOI21 U2166 (.OUT(n2482),
	.C(n2481),
	.B(n1433),
	.A(n1432));
   AOI21 U2167 (.OUT(n2483),
	.C(n2482),
	.B(\mult_19_3/ab[5][6] ),
	.A(\mult_19_3/ab[4][7] ));
   AOI21 U2168 (.OUT(n2484),
	.C(n2483),
	.B(n1435),
	.A(n1434));
   AOI21 U2169 (.OUT(n2485),
	.C(n2484),
	.B(\mult_19_3/ab[6][6] ),
	.A(\mult_19_3/ab[5][7] ));
   OAI21 U2170 (.OUT(n2486),
	.C(n2487),
	.B(\mult_19_3/ab[7][6] ),
	.A(\mult_19_3/ab[6][7] ));
   AOI21 U2171 (.OUT(n96),
	.C(n2488),
	.B(\mult_19_3/ab[7][6] ),
	.A(\mult_19_3/ab[6][7] ));
   AOI21 U2172 (.OUT(n1438),
	.C(n586),
	.B(n1395),
	.A(n2020));
   AOI21 U2173 (.OUT(n2489),
	.C(n609),
	.B(n1436),
	.A(n1439));
   OAI21 U2174 (.OUT(n2490),
	.C(n611),
	.B(n1440),
	.A(\mult_19_3/ab[7][5] ));
   AOI21 U2175 (.OUT(n98),
	.C(n2491),
	.B(\mult_19_3/ab[7][5] ),
	.A(n1440));
   OAI21 U2176 (.OUT(n2492),
	.C(n585),
	.B(n1397),
	.A(\mult_19_3/ab[6][4] ));
   inverter U2177 (.IN(n1442),
	.OUT(n2493));
   OAI21 U2178 (.OUT(n2494),
	.C(n608),
	.B(n2493),
	.A(\mult_19_3/ab[7][4] ));
   OAI21 U2179 (.OUT(n101),
	.C(n2494),
	.B(n2495),
	.A(n1442));
   OAI21 U2180 (.OUT(n2496),
	.C(n2497),
	.B(n1399),
	.A(\mult_19_3/ab[7][3] ));
   AOI21 U2181 (.OUT(n103),
	.C(n2498),
	.B(\mult_19_3/ab[7][3] ),
	.A(n1399));
   OAI21 U2182 (.OUT(n2499),
	.C(n2032),
	.B(\mult_19_2/ab[2][6] ),
	.A(\mult_19_2/ab[1][7] ));
   AOI21 U2183 (.OUT(n2500),
	.C(n2501),
	.B(\mult_19_2/ab[1][7] ),
	.A(\mult_19_2/ab[2][6] ));
   AOI21 U2184 (.OUT(n2502),
	.C(n2500),
	.B(n1481),
	.A(n1482));
   AOI21 U2185 (.OUT(n2503),
	.C(n2502),
	.B(\mult_19_2/ab[2][7] ),
	.A(\mult_19_2/ab[3][6] ));
   OAI21 U2186 (.OUT(n1472),
	.C(n618),
	.B(n2107),
	.A(\mult_19_2/ab[2][5] ));
   inverter U2187 (.IN(n1470),
	.OUT(n1484));
   OAI21 U2188 (.OUT(n1486),
	.C(n616),
	.B(n1470),
	.A(\mult_19_2/ab[3][5] ));
   OAI21 U2189 (.OUT(n2504),
	.C(n635),
	.B(n1483),
	.A(\mult_19_2/ab[4][5] ));
   inverter U2190 (.IN(n1495),
	.OUT(n1537));
   OAI21 U2191 (.OUT(n1463),
	.C(n619),
	.B(n2108),
	.A(\mult_19_2/ab[2][4] ));
   AOI21 U2192 (.OUT(n1475),
	.C(n620),
	.B(n2505),
	.A(n1460));
   AOI21 U2193 (.OUT(n1490),
	.C(n623),
	.B(n1474),
	.A(n1473));
   OAI21 U2194 (.OUT(n1498),
	.C(n634),
	.B(n2506),
	.A(\mult_19_2/ab[5][4] ));
   OAI21 U2195 (.OUT(n1456),
	.C(n625),
	.B(n2109),
	.A(\mult_19_2/ab[2][3] ));
   AOI21 U2196 (.OUT(n1465),
	.C(n626),
	.B(n2507),
	.A(n1453));
   inverter U2197 (.IN(n1464),
	.OUT(n2031));
   OAI21 U2198 (.OUT(n1478),
	.C(n632),
	.B(n2031),
	.A(\mult_19_2/ab[4][3] ));
   OAI21 U2199 (.OUT(n2508),
	.C(n622),
	.B(n1476),
	.A(\mult_19_2/ab[5][3] ));
   AOI21 U2200 (.OUT(n2509),
	.C(n638),
	.B(n1491),
	.A(n1500));
   OAI21 U2201 (.OUT(n2510),
	.C(n628),
	.B(n1446),
	.A(\mult_19_2/ab[2][2] ));
   AOI21 U2202 (.OUT(n2511),
	.C(n629),
	.B(n1445),
	.A(n1449));
   OAI21 U2203 (.OUT(n2512),
	.C(n649),
	.B(n1450),
	.A(\mult_19_2/ab[4][2] ));
   AOI21 U2204 (.OUT(n2513),
	.C(n631),
	.B(n1457),
	.A(n1466));
   OAI21 U2205 (.OUT(n2514),
	.C(n652),
	.B(n1467),
	.A(\mult_19_2/ab[6][2] ));
   inverter U2206 (.IN(n1479),
	.OUT(n2515));
   OAI21 U2207 (.OUT(n2516),
	.C(n637),
	.B(n2515),
	.A(\mult_19_2/ab[7][2] ));
   AOI21 U2208 (.OUT(n90),
	.C(n2517),
	.B(\mult_19_2/ab[7][2] ),
	.A(n2515));
   OAI21 U2209 (.OUT(n1505),
	.C(n645),
	.B(n2110),
	.A(\mult_19_2/ab[2][1] ));
   AOI21 U2210 (.OUT(n1508),
	.C(n646),
	.B(n2518),
	.A(n1506));
   inverter U2211 (.IN(n1507),
	.OUT(n2519));
   OAI21 U2212 (.OUT(n1511),
	.C(n658),
	.B(n2519),
	.A(\mult_19_2/ab[4][1] ));
   OAI21 U2213 (.OUT(n2520),
	.C(n648),
	.B(n1509),
	.A(\mult_19_2/ab[5][1] ));
   inverter U2214 (.IN(n1512),
	.OUT(n2521));
   OAI21 U2215 (.OUT(n1516),
	.C(n661),
	.B(n2521),
	.A(\mult_19_2/ab[6][1] ));
   OAI21 U2216 (.OUT(n2522),
	.C(n651),
	.B(n1515),
	.A(\mult_19_2/ab[7][1] ));
   AOI21 U2217 (.OUT(n92),
	.C(n2523),
	.B(\mult_19_2/ab[7][1] ),
	.A(n1515));
   OAI21 U2218 (.OUT(n2524),
	.C(n654),
	.B(n1519),
	.A(\mult_19_2/ab[2][0] ));
   AOI21 U2219 (.OUT(n2525),
	.C(n655),
	.B(n1518),
	.A(n1521));
   OAI21 U2220 (.OUT(n2526),
	.C(n1825),
	.B(n1522),
	.A(\mult_19_2/ab[4][0] ));
   AOI21 U2221 (.OUT(n2527),
	.C(n657),
	.B(n1524),
	.A(n1526));
   OAI21 U2222 (.OUT(n2528),
	.C(n1823),
	.B(n1527),
	.A(\mult_19_2/ab[6][0] ));
   inverter U2223 (.IN(n1529),
	.OUT(n2529));
   AOI21 U2224 (.OUT(n2530),
	.C(n660),
	.B(n1529),
	.A(n1531));
   AOI21 U2225 (.OUT(n94),
	.C(n2530),
	.B(\mult_19_2/ab[7][0] ),
	.A(n2529));
   AOI21 U2226 (.OUT(n2531),
	.C(n2503),
	.B(n1493),
	.A(n1494));
   AOI21 U2227 (.OUT(n2532),
	.C(n2531),
	.B(\mult_19_2/ab[3][7] ),
	.A(\mult_19_2/ab[4][6] ));
   AOI21 U2228 (.OUT(n2533),
	.C(n2532),
	.B(n1533),
	.A(n1532));
   AOI21 U2229 (.OUT(n2534),
	.C(n2533),
	.B(\mult_19_2/ab[5][6] ),
	.A(\mult_19_2/ab[4][7] ));
   AOI21 U2230 (.OUT(n2535),
	.C(n2534),
	.B(n1535),
	.A(n1534));
   AOI21 U2231 (.OUT(n2536),
	.C(n2535),
	.B(\mult_19_2/ab[6][6] ),
	.A(\mult_19_2/ab[5][7] ));
   OAI21 U2232 (.OUT(n2537),
	.C(n2538),
	.B(\mult_19_2/ab[7][6] ),
	.A(\mult_19_2/ab[6][7] ));
   AOI21 U2233 (.OUT(n81),
	.C(n2539),
	.B(\mult_19_2/ab[7][6] ),
	.A(\mult_19_2/ab[6][7] ));
   AOI21 U2234 (.OUT(n1538),
	.C(n641),
	.B(n1495),
	.A(n2036));
   AOI21 U2235 (.OUT(n2540),
	.C(n664),
	.B(n1536),
	.A(n1539));
   OAI21 U2236 (.OUT(n2541),
	.C(n666),
	.B(n1540),
	.A(\mult_19_2/ab[7][5] ));
   AOI21 U2237 (.OUT(n83),
	.C(n2542),
	.B(\mult_19_2/ab[7][5] ),
	.A(n1540));
   OAI21 U2238 (.OUT(n2543),
	.C(n640),
	.B(n1497),
	.A(\mult_19_2/ab[6][4] ));
   inverter U2239 (.IN(n1542),
	.OUT(n2544));
   OAI21 U2240 (.OUT(n2545),
	.C(n663),
	.B(n2544),
	.A(\mult_19_2/ab[7][4] ));
   OAI21 U2241 (.OUT(n86),
	.C(n2545),
	.B(n2546),
	.A(n1542));
   OAI21 U2242 (.OUT(n2547),
	.C(n2548),
	.B(n1499),
	.A(\mult_19_2/ab[7][3] ));
   AOI21 U2243 (.OUT(n88),
	.C(n2549),
	.B(\mult_19_2/ab[7][3] ),
	.A(n1499));
   OAI21 U2244 (.OUT(n2550),
	.C(n2048),
	.B(\mult_19/ab[2][6] ),
	.A(\mult_19/ab[1][7] ));
   AOI21 U2245 (.OUT(n2551),
	.C(n2552),
	.B(\mult_19/ab[1][7] ),
	.A(\mult_19/ab[2][6] ));
   AOI21 U2246 (.OUT(n2553),
	.C(n2551),
	.B(n1581),
	.A(n1582));
   AOI21 U2247 (.OUT(n2554),
	.C(n2553),
	.B(\mult_19/ab[2][7] ),
	.A(\mult_19/ab[3][6] ));
   OAI21 U2248 (.OUT(n1572),
	.C(n673),
	.B(n2103),
	.A(\mult_19/ab[2][5] ));
   inverter U2249 (.IN(n1570),
	.OUT(n1584));
   OAI21 U2250 (.OUT(n1586),
	.C(n671),
	.B(n1570),
	.A(\mult_19/ab[3][5] ));
   OAI21 U2251 (.OUT(n2555),
	.C(n690),
	.B(n1583),
	.A(\mult_19/ab[4][5] ));
   inverter U2252 (.IN(n1595),
	.OUT(n1637));
   OAI21 U2253 (.OUT(n1563),
	.C(n674),
	.B(n2104),
	.A(\mult_19/ab[2][4] ));
   AOI21 U2254 (.OUT(n1575),
	.C(n675),
	.B(n2556),
	.A(n1560));
   AOI21 U2255 (.OUT(n1590),
	.C(n678),
	.B(n1574),
	.A(n1573));
   OAI21 U2256 (.OUT(n1598),
	.C(n689),
	.B(n2557),
	.A(\mult_19/ab[5][4] ));
   OAI21 U2257 (.OUT(n1556),
	.C(n680),
	.B(n2105),
	.A(\mult_19/ab[2][3] ));
   AOI21 U2258 (.OUT(n1565),
	.C(n681),
	.B(n2558),
	.A(n1553));
   inverter U2259 (.IN(n1564),
	.OUT(n2047));
   OAI21 U2260 (.OUT(n1578),
	.C(n687),
	.B(n2047),
	.A(\mult_19/ab[4][3] ));
   OAI21 U2261 (.OUT(n2559),
	.C(n677),
	.B(n1576),
	.A(\mult_19/ab[5][3] ));
   AOI21 U2262 (.OUT(n2560),
	.C(n693),
	.B(n1591),
	.A(n1600));
   OAI21 U2263 (.OUT(n2561),
	.C(n683),
	.B(n1546),
	.A(\mult_19/ab[2][2] ));
   AOI21 U2264 (.OUT(n2562),
	.C(n684),
	.B(n1545),
	.A(n1549));
   OAI21 U2265 (.OUT(n2563),
	.C(n704),
	.B(n1550),
	.A(\mult_19/ab[4][2] ));
   AOI21 U2266 (.OUT(n2564),
	.C(n686),
	.B(n1557),
	.A(n1566));
   OAI21 U2267 (.OUT(n2565),
	.C(n707),
	.B(n1567),
	.A(\mult_19/ab[6][2] ));
   inverter U2268 (.IN(n1579),
	.OUT(n2566));
   OAI21 U2269 (.OUT(n2567),
	.C(n692),
	.B(n2566),
	.A(\mult_19/ab[7][2] ));
   AOI21 U2270 (.OUT(n75),
	.C(n2568),
	.B(\mult_19/ab[7][2] ),
	.A(n2566));
   OAI21 U2271 (.OUT(n1605),
	.C(n700),
	.B(n2106),
	.A(\mult_19/ab[2][1] ));
   AOI21 U2272 (.OUT(n1608),
	.C(n701),
	.B(n2569),
	.A(n1606));
   inverter U2273 (.IN(n1607),
	.OUT(n2570));
   OAI21 U2274 (.OUT(n1611),
	.C(n713),
	.B(n2570),
	.A(\mult_19/ab[4][1] ));
   OAI21 U2275 (.OUT(n2571),
	.C(n703),
	.B(n1609),
	.A(\mult_19/ab[5][1] ));
   inverter U2276 (.IN(n1612),
	.OUT(n2572));
   OAI21 U2277 (.OUT(n1616),
	.C(n716),
	.B(n2572),
	.A(\mult_19/ab[6][1] ));
   OAI21 U2278 (.OUT(n2573),
	.C(n706),
	.B(n1615),
	.A(\mult_19/ab[7][1] ));
   AOI21 U2279 (.OUT(n77),
	.C(n2574),
	.B(\mult_19/ab[7][1] ),
	.A(n1615));
   OAI21 U2280 (.OUT(n2575),
	.C(n709),
	.B(n1619),
	.A(\mult_19/ab[2][0] ));
   AOI21 U2281 (.OUT(n2576),
	.C(n710),
	.B(n1618),
	.A(n1621));
   OAI21 U2282 (.OUT(n2577),
	.C(n1830),
	.B(n1622),
	.A(\mult_19/ab[4][0] ));
   AOI21 U2283 (.OUT(n2578),
	.C(n712),
	.B(n1624),
	.A(n1626));
   OAI21 U2284 (.OUT(n2579),
	.C(n1828),
	.B(n1627),
	.A(\mult_19/ab[6][0] ));
   inverter U2285 (.IN(n1629),
	.OUT(n2580));
   AOI21 U2286 (.OUT(n2581),
	.C(n715),
	.B(n1629),
	.A(n1631));
   AOI21 U2287 (.OUT(n79),
	.C(n2581),
	.B(\mult_19/ab[7][0] ),
	.A(n2580));
   AOI21 U2288 (.OUT(n2582),
	.C(n2554),
	.B(n1593),
	.A(n1594));
   AOI21 U2289 (.OUT(n2583),
	.C(n2582),
	.B(\mult_19/ab[3][7] ),
	.A(\mult_19/ab[4][6] ));
   AOI21 U2290 (.OUT(n2584),
	.C(n2583),
	.B(n1633),
	.A(n1632));
   AOI21 U2291 (.OUT(n2585),
	.C(n2584),
	.B(\mult_19/ab[5][6] ),
	.A(\mult_19/ab[4][7] ));
   AOI21 U2292 (.OUT(n2586),
	.C(n2585),
	.B(n1635),
	.A(n1634));
   AOI21 U2293 (.OUT(n2587),
	.C(n2586),
	.B(\mult_19/ab[6][6] ),
	.A(\mult_19/ab[5][7] ));
   OAI21 U2294 (.OUT(n2588),
	.C(n2589),
	.B(\mult_19/ab[7][6] ),
	.A(\mult_19/ab[6][7] ));
   AOI21 U2295 (.OUT(n66),
	.C(n2590),
	.B(\mult_19/ab[7][6] ),
	.A(\mult_19/ab[6][7] ));
   AOI21 U2296 (.OUT(n1638),
	.C(n696),
	.B(n1595),
	.A(n2052));
   AOI21 U2297 (.OUT(n2591),
	.C(n719),
	.B(n1636),
	.A(n1639));
   OAI21 U2298 (.OUT(n2592),
	.C(n721),
	.B(n1640),
	.A(\mult_19/ab[7][5] ));
   AOI21 U2299 (.OUT(n68),
	.C(n2593),
	.B(\mult_19/ab[7][5] ),
	.A(n1640));
   OAI21 U2300 (.OUT(n2594),
	.C(n695),
	.B(n1597),
	.A(\mult_19/ab[6][4] ));
   inverter U2301 (.IN(n1642),
	.OUT(n2595));
   OAI21 U2302 (.OUT(n2596),
	.C(n718),
	.B(n2595),
	.A(\mult_19/ab[7][4] ));
   OAI21 U2303 (.OUT(n71),
	.C(n2596),
	.B(n2597),
	.A(n1642));
   OAI21 U2304 (.OUT(n2598),
	.C(n2599),
	.B(n1599),
	.A(\mult_19/ab[7][3] ));
   AOI21 U2305 (.OUT(n73),
	.C(n2600),
	.B(\mult_19/ab[7][3] ),
	.A(n1599));
   OAI21 U2306 (.OUT(n2601),
	.C(n727),
	.B(n726),
	.A(n2111));
   OAI21 U2307 (.OUT(n2602),
	.C(n2601),
	.B(n1644),
	.A(n2603));
   OAI21 U2308 (.OUT(n2604),
	.C(n2602),
	.B(N3),
	.A(N19));
   AOI21 U2309 (.OUT(n2605),
	.C(n2606),
	.B(N3),
	.A(N19));
   OAI21 U2310 (.OUT(n2607),
	.C(n2608),
	.B(N4),
	.A(N20));
   AOI21 U2311 (.OUT(n2609),
	.C(n2610),
	.B(N4),
	.A(N20));
   OAI21 U2312 (.OUT(n2611),
	.C(n2612),
	.B(N5),
	.A(N21));
   AOI21 U2313 (.OUT(n2613),
	.C(n2614),
	.B(N5),
	.A(N21));
   OAI21 U2314 (.OUT(n2615),
	.C(n2616),
	.B(N6),
	.A(N22));
   AOI21 U2315 (.OUT(n2617),
	.C(n2618),
	.B(N6),
	.A(N22));
   OAI21 U2316 (.OUT(n2619),
	.C(n2620),
	.B(N7),
	.A(N23));
   AOI21 U2317 (.OUT(n2621),
	.C(n2622),
	.B(N7),
	.A(N23));
   OAI21 U2318 (.OUT(n2623),
	.C(n2624),
	.B(N8),
	.A(N24));
   AOI21 U2319 (.OUT(n2625),
	.C(n2626),
	.B(N8),
	.A(N24));
   OAI21 U2320 (.OUT(n2627),
	.C(n2628),
	.B(N9),
	.A(N25));
   AOI21 U2321 (.OUT(n2629),
	.C(n2630),
	.B(N9),
	.A(N25));
   OAI21 U2322 (.OUT(n2631),
	.C(n2632),
	.B(N10),
	.A(N26));
   AOI21 U2323 (.OUT(n2633),
	.C(n2634),
	.B(N10),
	.A(N26));
   OAI21 U2324 (.OUT(n2635),
	.C(n2636),
	.B(N11),
	.A(N27));
   AOI21 U2325 (.OUT(n2637),
	.C(n2638),
	.B(N11),
	.A(N27));
   OAI21 U2326 (.OUT(n2639),
	.C(n2640),
	.B(N12),
	.A(N28));
   AOI21 U2327 (.OUT(n2641),
	.C(n2642),
	.B(N12),
	.A(N28));
   OAI21 U2328 (.OUT(n2643),
	.C(n2644),
	.B(N13),
	.A(N29));
   AOI21 U2329 (.OUT(n2645),
	.C(n2646),
	.B(N13),
	.A(N29));
   OAI21 U2330 (.OUT(n2647),
	.C(n2648),
	.B(N14),
	.A(N30));
   AOI21 U2331 (.OUT(n2649),
	.C(n2650),
	.B(N14),
	.A(N30));
   OAI21 U2332 (.OUT(n1648),
	.C(n730),
	.B(n729),
	.A(n2074));
   OAI21 U2333 (.OUT(n2651),
	.C(n1858),
	.B(n1646),
	.A(N51));
   AOI21 U2334 (.OUT(n2652),
	.C(n1856),
	.B(n1649),
	.A(n1651));
   AOI21 U2335 (.OUT(n1656),
	.C(n1854),
	.B(n2653),
	.A(n1654));
   AOI21 U2336 (.OUT(n1660),
	.C(n1852),
	.B(n1655),
	.A(n1657));
   AOI21 U2337 (.OUT(n1664),
	.C(n1850),
	.B(n1658),
	.A(n1661));
   AOI21 U2338 (.OUT(n1668),
	.C(n1848),
	.B(n1662),
	.A(n1665));
   AOI21 U2339 (.OUT(n1672),
	.C(n1846),
	.B(n1666),
	.A(n1669));
   AOI21 U2340 (.OUT(n1676),
	.C(n1844),
	.B(n1670),
	.A(n1673));
   AOI21 U2341 (.OUT(n1680),
	.C(n1842),
	.B(n1674),
	.A(n1677));
   AOI21 U2342 (.OUT(n1684),
	.C(n1840),
	.B(n1678),
	.A(n1681));
   AOI21 U2343 (.OUT(n1688),
	.C(n1838),
	.B(n1682),
	.A(n1685));
   AOI21 U2344 (.OUT(n1691),
	.C(n1836),
	.B(n1686),
	.A(n1689));
   inverter U2345 (.IN(n206),
	.OUT(n210));
   OAI21 U2346 (.OUT(n2654),
	.C(n733),
	.B(n732),
	.A(n2137));
   OAI21 U2347 (.OUT(n2655),
	.C(n2654),
	.B(n1692),
	.A(n2656));
   OAI21 U2348 (.OUT(n2657),
	.C(n2655),
	.B(N163),
	.A(N179));
   AOI21 U2349 (.OUT(n2658),
	.C(n2659),
	.B(N163),
	.A(N179));
   OAI21 U2350 (.OUT(n2660),
	.C(n2661),
	.B(N164),
	.A(N180));
   AOI21 U2351 (.OUT(n2662),
	.C(n2663),
	.B(N164),
	.A(N180));
   OAI21 U2352 (.OUT(n2664),
	.C(n2665),
	.B(N165),
	.A(N181));
   AOI21 U2353 (.OUT(n2666),
	.C(n2667),
	.B(N165),
	.A(N181));
   OAI21 U2354 (.OUT(n2668),
	.C(n2669),
	.B(N166),
	.A(N182));
   AOI21 U2355 (.OUT(n2670),
	.C(n2671),
	.B(N166),
	.A(N182));
   OAI21 U2356 (.OUT(n2672),
	.C(n2673),
	.B(N167),
	.A(N183));
   AOI21 U2357 (.OUT(n2674),
	.C(n2675),
	.B(N167),
	.A(N183));
   OAI21 U2358 (.OUT(n2676),
	.C(n2677),
	.B(N168),
	.A(N184));
   AOI21 U2359 (.OUT(n2678),
	.C(n2679),
	.B(N168),
	.A(N184));
   OAI21 U2360 (.OUT(n2680),
	.C(n2681),
	.B(N169),
	.A(N185));
   AOI21 U2361 (.OUT(n2682),
	.C(n2683),
	.B(N169),
	.A(N185));
   OAI21 U2362 (.OUT(n2684),
	.C(n2685),
	.B(N170),
	.A(N186));
   AOI21 U2363 (.OUT(n2686),
	.C(n2687),
	.B(N170),
	.A(N186));
   OAI21 U2364 (.OUT(n2688),
	.C(n2689),
	.B(N171),
	.A(N187));
   AOI21 U2365 (.OUT(n2690),
	.C(n2691),
	.B(N171),
	.A(N187));
   OAI21 U2366 (.OUT(n2692),
	.C(n2693),
	.B(N172),
	.A(N188));
   AOI21 U2367 (.OUT(n2694),
	.C(n2695),
	.B(N172),
	.A(N188));
   OAI21 U2368 (.OUT(n2696),
	.C(n2697),
	.B(N173),
	.A(N189));
   AOI21 U2369 (.OUT(n2698),
	.C(n2699),
	.B(N173),
	.A(N189));
   OAI21 U2370 (.OUT(n2700),
	.C(n2701),
	.B(N174),
	.A(N190));
   AOI21 U2371 (.OUT(n2702),
	.C(n2703),
	.B(N174),
	.A(N190));
   OAI21 U2372 (.OUT(n1696),
	.C(n736),
	.B(n735),
	.A(n2088));
   OAI21 U2373 (.OUT(n2704),
	.C(n1886),
	.B(n1694),
	.A(N211));
   AOI21 U2374 (.OUT(n2705),
	.C(n1884),
	.B(n1697),
	.A(n1699));
   AOI21 U2375 (.OUT(n1704),
	.C(n1882),
	.B(n2706),
	.A(n1702));
   AOI21 U2376 (.OUT(n1708),
	.C(n1880),
	.B(n1703),
	.A(n1705));
   AOI21 U2377 (.OUT(n1712),
	.C(n1878),
	.B(n1706),
	.A(n1709));
   AOI21 U2378 (.OUT(n1716),
	.C(n1876),
	.B(n1710),
	.A(n1713));
   AOI21 U2379 (.OUT(n1720),
	.C(n1874),
	.B(n1714),
	.A(n1717));
   AOI21 U2380 (.OUT(n1724),
	.C(n1872),
	.B(n1718),
	.A(n1721));
   AOI21 U2381 (.OUT(n1728),
	.C(n1870),
	.B(n1722),
	.A(n1725));
   AOI21 U2382 (.OUT(n1732),
	.C(n1868),
	.B(n1726),
	.A(n1729));
   AOI21 U2383 (.OUT(n1736),
	.C(n1866),
	.B(n1730),
	.A(n1733));
   AOI21 U2384 (.OUT(n1739),
	.C(n1864),
	.B(n1734),
	.A(n1737));
   inverter U2385 (.IN(n216),
	.OUT(n220));
   OAI21 U2386 (.OUT(n2707),
	.C(n739),
	.B(n738),
	.A(n2124));
   OAI21 U2387 (.OUT(n2708),
	.C(n2707),
	.B(n1740),
	.A(n2709));
   OAI21 U2388 (.OUT(n2710),
	.C(n2708),
	.B(N83),
	.A(N99));
   AOI21 U2389 (.OUT(n2711),
	.C(n2712),
	.B(N83),
	.A(N99));
   OAI21 U2390 (.OUT(n2713),
	.C(n2714),
	.B(N84),
	.A(N100));
   AOI21 U2391 (.OUT(n2715),
	.C(n2716),
	.B(N84),
	.A(N100));
   OAI21 U2392 (.OUT(n2717),
	.C(n2718),
	.B(N85),
	.A(N101));
   AOI21 U2393 (.OUT(n2719),
	.C(n2720),
	.B(N85),
	.A(N101));
   OAI21 U2394 (.OUT(n2721),
	.C(n2722),
	.B(N86),
	.A(N102));
   AOI21 U2395 (.OUT(n2723),
	.C(n2724),
	.B(N86),
	.A(N102));
   OAI21 U2396 (.OUT(n2725),
	.C(n2726),
	.B(N87),
	.A(N103));
   AOI21 U2397 (.OUT(n2727),
	.C(n2728),
	.B(N87),
	.A(N103));
   OAI21 U2398 (.OUT(n2729),
	.C(n2730),
	.B(N88),
	.A(N104));
   AOI21 U2399 (.OUT(n2731),
	.C(n2732),
	.B(N88),
	.A(N104));
   OAI21 U2400 (.OUT(n2733),
	.C(n2734),
	.B(N89),
	.A(N105));
   AOI21 U2401 (.OUT(n2735),
	.C(n2736),
	.B(N89),
	.A(N105));
   OAI21 U2402 (.OUT(n2737),
	.C(n2738),
	.B(N90),
	.A(N106));
   AOI21 U2403 (.OUT(n2739),
	.C(n2740),
	.B(N90),
	.A(N106));
   OAI21 U2404 (.OUT(n2741),
	.C(n2742),
	.B(N91),
	.A(N107));
   AOI21 U2405 (.OUT(n2743),
	.C(n2744),
	.B(N91),
	.A(N107));
   OAI21 U2406 (.OUT(n2745),
	.C(n2746),
	.B(N92),
	.A(N108));
   AOI21 U2407 (.OUT(n2747),
	.C(n2748),
	.B(N92),
	.A(N108));
   OAI21 U2408 (.OUT(n2749),
	.C(n2750),
	.B(N93),
	.A(N109));
   AOI21 U2409 (.OUT(n2751),
	.C(n2752),
	.B(N93),
	.A(N109));
   OAI21 U2410 (.OUT(n2753),
	.C(n2754),
	.B(N94),
	.A(N110));
   AOI21 U2411 (.OUT(n2755),
	.C(n2756),
	.B(N94),
	.A(N110));
   OAI21 U2412 (.OUT(n1744),
	.C(n742),
	.B(n741),
	.A(n2102));
   OAI21 U2413 (.OUT(n2757),
	.C(n1914),
	.B(n1742),
	.A(N131));
   AOI21 U2414 (.OUT(n2758),
	.C(n1912),
	.B(n1745),
	.A(n1747));
   AOI21 U2415 (.OUT(n1752),
	.C(n1910),
	.B(n2759),
	.A(n1750));
   AOI21 U2416 (.OUT(n1756),
	.C(n1908),
	.B(n1751),
	.A(n1753));
   AOI21 U2417 (.OUT(n1760),
	.C(n1906),
	.B(n1754),
	.A(n1757));
   AOI21 U2418 (.OUT(n1764),
	.C(n1904),
	.B(n1758),
	.A(n1761));
   AOI21 U2419 (.OUT(n1768),
	.C(n1902),
	.B(n1762),
	.A(n1765));
   AOI21 U2420 (.OUT(n1772),
	.C(n1900),
	.B(n1766),
	.A(n1769));
   AOI21 U2421 (.OUT(n1776),
	.C(n1898),
	.B(n1770),
	.A(n1773));
   AOI21 U2422 (.OUT(n1780),
	.C(n1896),
	.B(n1774),
	.A(n1777));
   AOI21 U2423 (.OUT(n1784),
	.C(n1894),
	.B(n1778),
	.A(n1781));
   AOI21 U2424 (.OUT(n1787),
	.C(n1892),
	.B(n1782),
	.A(n1785));
   inverter U2425 (.IN(n226),
	.OUT(n230));
   XOR2 U2426 (.A(n241),
	.B(n1917),
	.OUT(n264));
   XOR2 U2427 (.A(n235),
	.B(n1918),
	.OUT(n247));
   XOR2 U2428 (.A(n231),
	.B(n1921),
	.OUT(n238));
   XOR2 U2429 (.A(n237),
	.B(n1922),
	.OUT(n267));
   XOR2 U2430 (.A(n2760),
	.B(n2143),
	.OUT(n250));
   XOR2 U2431 (.A(n249),
	.B(n1923),
	.OUT(n253));
   XOR2 U2432 (.A(n2761),
	.B(n2146),
	.OUT(n256));
   XOR2 U2433 (.A(n255),
	.B(n1925),
	.OUT(n2191));
   XOR2 U2434 (.A(n244),
	.B(n1926),
	.OUT(n273));
   XOR2 U2435 (.A(n246),
	.B(n1927),
	.OUT(n276));
   XOR2 U2436 (.A(n252),
	.B(n1928),
	.OUT(n198));
   XOR2 U2437 (.A(n261),
	.B(n1929),
	.OUT(n1790));
   XOR2 U2438 (.A(n263),
	.B(n1930),
	.OUT(n1788));
   XOR2 U2439 (.A(n266),
	.B(n1931),
	.OUT(n2762));
   XOR2 U2440 (.A(n2763),
	.B(n2175),
	.OUT(n279));
   XOR2 U2441 (.A(n2764),
	.B(n2177),
	.OUT(n281));
   XOR2 U2442 (.A(n2765),
	.B(n2179),
	.OUT(n189));
   XOR2 U2443 (.A(n278),
	.B(n1932),
	.OUT(n194));
   XOR2 U2444 (.A(n296),
	.B(n1933),
	.OUT(n319));
   XOR2 U2445 (.A(n290),
	.B(n1934),
	.OUT(n302));
   XOR2 U2446 (.A(n286),
	.B(n1937),
	.OUT(n293));
   XOR2 U2447 (.A(n292),
	.B(n1938),
	.OUT(n322));
   XOR2 U2448 (.A(n2766),
	.B(n2194),
	.OUT(n305));
   XOR2 U2449 (.A(n304),
	.B(n1939),
	.OUT(n308));
   XOR2 U2450 (.A(n2767),
	.B(n2197),
	.OUT(n311));
   XOR2 U2451 (.A(n310),
	.B(n1941),
	.OUT(n2242));
   XOR2 U2452 (.A(n299),
	.B(n1942),
	.OUT(n328));
   XOR2 U2453 (.A(n301),
	.B(n1943),
	.OUT(n331));
   XOR2 U2454 (.A(n307),
	.B(n1944),
	.OUT(n183));
   XOR2 U2455 (.A(n316),
	.B(n1945),
	.OUT(n1795));
   XOR2 U2456 (.A(n318),
	.B(n1946),
	.OUT(n1793));
   XOR2 U2457 (.A(n321),
	.B(n1947),
	.OUT(n2768));
   XOR2 U2458 (.A(n2769),
	.B(n2226),
	.OUT(n334));
   XOR2 U2459 (.A(n2770),
	.B(n2228),
	.OUT(n336));
   XOR2 U2460 (.A(n2771),
	.B(n2230),
	.OUT(n174));
   XOR2 U2461 (.A(n333),
	.B(n1948),
	.OUT(n179));
   XOR2 U2462 (.A(n351),
	.B(n1949),
	.OUT(n374));
   XOR2 U2463 (.A(n345),
	.B(n1950),
	.OUT(n357));
   XOR2 U2464 (.A(n341),
	.B(n1953),
	.OUT(n348));
   XOR2 U2465 (.A(n347),
	.B(n1954),
	.OUT(n377));
   XOR2 U2466 (.A(n2772),
	.B(n2245),
	.OUT(n360));
   XOR2 U2467 (.A(n359),
	.B(n1955),
	.OUT(n363));
   XOR2 U2468 (.A(n2773),
	.B(n2248),
	.OUT(n366));
   XOR2 U2469 (.A(n365),
	.B(n1957),
	.OUT(n2293));
   XOR2 U2470 (.A(n354),
	.B(n1958),
	.OUT(n383));
   XOR2 U2471 (.A(n356),
	.B(n1959),
	.OUT(n386));
   XOR2 U2472 (.A(n362),
	.B(n1960),
	.OUT(n168));
   XOR2 U2473 (.A(n371),
	.B(n1961),
	.OUT(n1800));
   XOR2 U2474 (.A(n373),
	.B(n1962),
	.OUT(n1798));
   XOR2 U2475 (.A(n376),
	.B(n1963),
	.OUT(n2774));
   XOR2 U2476 (.A(n2775),
	.B(n2277),
	.OUT(n389));
   XOR2 U2477 (.A(n2776),
	.B(n2279),
	.OUT(n391));
   XOR2 U2478 (.A(n2777),
	.B(n2281),
	.OUT(n159));
   XOR2 U2479 (.A(n388),
	.B(n1964),
	.OUT(n164));
   XOR2 U2480 (.A(n406),
	.B(n1965),
	.OUT(n429));
   XOR2 U2481 (.A(n400),
	.B(n1966),
	.OUT(n412));
   XOR2 U2482 (.A(n396),
	.B(n1969),
	.OUT(n403));
   XOR2 U2483 (.A(n402),
	.B(n1970),
	.OUT(n432));
   XOR2 U2484 (.A(n2778),
	.B(n2296),
	.OUT(n415));
   XOR2 U2485 (.A(n414),
	.B(n1971),
	.OUT(n418));
   XOR2 U2486 (.A(n2779),
	.B(n2299),
	.OUT(n421));
   XOR2 U2487 (.A(n420),
	.B(n1973),
	.OUT(n2344));
   XOR2 U2488 (.A(n409),
	.B(n1974),
	.OUT(n438));
   XOR2 U2489 (.A(n411),
	.B(n1975),
	.OUT(n441));
   XOR2 U2490 (.A(n417),
	.B(n1976),
	.OUT(n153));
   XOR2 U2491 (.A(n426),
	.B(n1977),
	.OUT(n1805));
   XOR2 U2492 (.A(n428),
	.B(n1978),
	.OUT(n1803));
   XOR2 U2493 (.A(n431),
	.B(n1979),
	.OUT(n2780));
   XOR2 U2494 (.A(n2781),
	.B(n2328),
	.OUT(n444));
   XOR2 U2495 (.A(n2782),
	.B(n2330),
	.OUT(n446));
   XOR2 U2496 (.A(n2783),
	.B(n2332),
	.OUT(n144));
   XOR2 U2497 (.A(n443),
	.B(n1980),
	.OUT(n149));
   XOR2 U2498 (.A(n461),
	.B(n1981),
	.OUT(n484));
   XOR2 U2499 (.A(n455),
	.B(n1982),
	.OUT(n467));
   XOR2 U2500 (.A(n451),
	.B(n1985),
	.OUT(n458));
   XOR2 U2501 (.A(n457),
	.B(n1986),
	.OUT(n487));
   XOR2 U2502 (.A(n2784),
	.B(n2347),
	.OUT(n470));
   XOR2 U2503 (.A(n469),
	.B(n1987),
	.OUT(n473));
   XOR2 U2504 (.A(n2785),
	.B(n2350),
	.OUT(n476));
   XOR2 U2505 (.A(n475),
	.B(n1989),
	.OUT(n2395));
   XOR2 U2506 (.A(n464),
	.B(n1990),
	.OUT(n493));
   XOR2 U2507 (.A(n466),
	.B(n1991),
	.OUT(n496));
   XOR2 U2508 (.A(n472),
	.B(n1992),
	.OUT(n138));
   XOR2 U2509 (.A(n481),
	.B(n1993),
	.OUT(n1810));
   XOR2 U2510 (.A(n483),
	.B(n1994),
	.OUT(n1808));
   XOR2 U2511 (.A(n486),
	.B(n1995),
	.OUT(n2786));
   XOR2 U2512 (.A(n2787),
	.B(n2379),
	.OUT(n499));
   XOR2 U2513 (.A(n2788),
	.B(n2381),
	.OUT(n501));
   XOR2 U2514 (.A(n2789),
	.B(n2383),
	.OUT(n129));
   XOR2 U2515 (.A(n498),
	.B(n1996),
	.OUT(n134));
   XOR2 U2516 (.A(n516),
	.B(n1997),
	.OUT(n539));
   XOR2 U2517 (.A(n510),
	.B(n1998),
	.OUT(n522));
   XOR2 U2518 (.A(n506),
	.B(n2001),
	.OUT(n513));
   XOR2 U2519 (.A(n512),
	.B(n2002),
	.OUT(n542));
   XOR2 U2520 (.A(n2790),
	.B(n2398),
	.OUT(n525));
   XOR2 U2521 (.A(n524),
	.B(n2003),
	.OUT(n528));
   XOR2 U2522 (.A(n2791),
	.B(n2401),
	.OUT(n531));
   XOR2 U2523 (.A(n530),
	.B(n2005),
	.OUT(n2446));
   XOR2 U2524 (.A(n519),
	.B(n2006),
	.OUT(n548));
   XOR2 U2525 (.A(n521),
	.B(n2007),
	.OUT(n551));
   XOR2 U2526 (.A(n527),
	.B(n2008),
	.OUT(n123));
   XOR2 U2527 (.A(n536),
	.B(n2009),
	.OUT(n1815));
   XOR2 U2528 (.A(n538),
	.B(n2010),
	.OUT(n1813));
   XOR2 U2529 (.A(n541),
	.B(n2011),
	.OUT(n2792));
   XOR2 U2530 (.A(n2793),
	.B(n2430),
	.OUT(n554));
   XOR2 U2531 (.A(n2794),
	.B(n2432),
	.OUT(n556));
   XOR2 U2532 (.A(n2795),
	.B(n2434),
	.OUT(n114));
   XOR2 U2533 (.A(n553),
	.B(n2012),
	.OUT(n119));
   XOR2 U2534 (.A(n571),
	.B(n2013),
	.OUT(n594));
   XOR2 U2535 (.A(n565),
	.B(n2014),
	.OUT(n577));
   XOR2 U2536 (.A(n561),
	.B(n2017),
	.OUT(n568));
   XOR2 U2537 (.A(n567),
	.B(n2018),
	.OUT(n597));
   XOR2 U2538 (.A(n2796),
	.B(n2449),
	.OUT(n580));
   XOR2 U2539 (.A(n579),
	.B(n2019),
	.OUT(n583));
   XOR2 U2540 (.A(n2797),
	.B(n2452),
	.OUT(n586));
   XOR2 U2541 (.A(n585),
	.B(n2021),
	.OUT(n2497));
   XOR2 U2542 (.A(n574),
	.B(n2022),
	.OUT(n603));
   XOR2 U2543 (.A(n576),
	.B(n2023),
	.OUT(n606));
   XOR2 U2544 (.A(n582),
	.B(n2024),
	.OUT(n108));
   XOR2 U2545 (.A(n591),
	.B(n2025),
	.OUT(n1820));
   XOR2 U2546 (.A(n593),
	.B(n2026),
	.OUT(n1818));
   XOR2 U2547 (.A(n596),
	.B(n2027),
	.OUT(n2798));
   XOR2 U2548 (.A(n2799),
	.B(n2481),
	.OUT(n609));
   XOR2 U2549 (.A(n2800),
	.B(n2483),
	.OUT(n611));
   XOR2 U2550 (.A(n2801),
	.B(n2485),
	.OUT(n99));
   XOR2 U2551 (.A(n608),
	.B(n2028),
	.OUT(n104));
   XOR2 U2552 (.A(n626),
	.B(n2029),
	.OUT(n649));
   XOR2 U2553 (.A(n620),
	.B(n2030),
	.OUT(n632));
   XOR2 U2554 (.A(n616),
	.B(n2033),
	.OUT(n623));
   XOR2 U2555 (.A(n622),
	.B(n2034),
	.OUT(n652));
   XOR2 U2556 (.A(n2802),
	.B(n2500),
	.OUT(n635));
   XOR2 U2557 (.A(n634),
	.B(n2035),
	.OUT(n638));
   XOR2 U2558 (.A(n2803),
	.B(n2503),
	.OUT(n641));
   XOR2 U2559 (.A(n640),
	.B(n2037),
	.OUT(n2548));
   XOR2 U2560 (.A(n629),
	.B(n2038),
	.OUT(n658));
   XOR2 U2561 (.A(n631),
	.B(n2039),
	.OUT(n661));
   XOR2 U2562 (.A(n637),
	.B(n2040),
	.OUT(n93));
   XOR2 U2563 (.A(n646),
	.B(n2041),
	.OUT(n1825));
   XOR2 U2564 (.A(n648),
	.B(n2042),
	.OUT(n1823));
   XOR2 U2565 (.A(n651),
	.B(n2043),
	.OUT(n2804));
   XOR2 U2566 (.A(n2805),
	.B(n2532),
	.OUT(n664));
   XOR2 U2567 (.A(n2806),
	.B(n2534),
	.OUT(n666));
   XOR2 U2568 (.A(n2807),
	.B(n2536),
	.OUT(n84));
   XOR2 U2569 (.A(n663),
	.B(n2044),
	.OUT(n89));
   XOR2 U2570 (.A(n681),
	.B(n2045),
	.OUT(n704));
   XOR2 U2571 (.A(n675),
	.B(n2046),
	.OUT(n687));
   XOR2 U2572 (.A(n671),
	.B(n2049),
	.OUT(n678));
   XOR2 U2573 (.A(n677),
	.B(n2050),
	.OUT(n707));
   XOR2 U2574 (.A(n2808),
	.B(n2551),
	.OUT(n690));
   XOR2 U2575 (.A(n689),
	.B(n2051),
	.OUT(n693));
   XOR2 U2576 (.A(n2809),
	.B(n2554),
	.OUT(n696));
   XOR2 U2577 (.A(n695),
	.B(n2053),
	.OUT(n2599));
   XOR2 U2578 (.A(n684),
	.B(n2054),
	.OUT(n713));
   XOR2 U2579 (.A(n686),
	.B(n2055),
	.OUT(n716));
   XOR2 U2580 (.A(n692),
	.B(n2056),
	.OUT(n78));
   XOR2 U2581 (.A(n701),
	.B(n2057),
	.OUT(n1830));
   XOR2 U2582 (.A(n703),
	.B(n2058),
	.OUT(n1828));
   XOR2 U2583 (.A(n706),
	.B(n2059),
	.OUT(n2810));
   XOR2 U2584 (.A(n2811),
	.B(n2583),
	.OUT(n719));
   XOR2 U2585 (.A(n2812),
	.B(n2585),
	.OUT(n721));
   XOR2 U2586 (.A(n2813),
	.B(n2587),
	.OUT(n69));
   XOR2 U2587 (.A(n718),
	.B(n2060),
	.OUT(n74));
   inverter U2588 (.IN(n729),
	.OUT(n1647));
   inverter U2589 (.IN(n726),
	.OUT(n2603));
   XOR2 U2590 (.A(n2602),
	.B(n2061),
	.OUT(n1858));
   XOR2 U2591 (.A(n2605),
	.B(n2062),
	.OUT(n1856));
   XOR2 U2592 (.A(n2609),
	.B(n2063),
	.OUT(n1854));
   XOR2 U2593 (.A(n2613),
	.B(n2064),
	.OUT(n1852));
   XOR2 U2594 (.A(n2617),
	.B(n2065),
	.OUT(n1850));
   XOR2 U2595 (.A(n2621),
	.B(n2066),
	.OUT(n1848));
   XOR2 U2596 (.A(n2625),
	.B(n2067),
	.OUT(n1846));
   XOR2 U2597 (.A(n2629),
	.B(n2068),
	.OUT(n1844));
   XOR2 U2598 (.A(n2633),
	.B(n2069),
	.OUT(n1842));
   XOR2 U2599 (.A(n2637),
	.B(n2070),
	.OUT(n1840));
   XOR2 U2600 (.A(n2641),
	.B(n2071),
	.OUT(n1838));
   XOR2 U2601 (.A(n2645),
	.B(n2072),
	.OUT(n1836));
   XOR2 U2602 (.A(n2814),
	.B(n2649),
	.OUT(n208));
   inverter U2603 (.IN(n735),
	.OUT(n1695));
   inverter U2604 (.IN(n732),
	.OUT(n2656));
   XOR2 U2605 (.A(n2655),
	.B(n2075),
	.OUT(n1886));
   XOR2 U2606 (.A(n2658),
	.B(n2076),
	.OUT(n1884));
   XOR2 U2607 (.A(n2662),
	.B(n2077),
	.OUT(n1882));
   XOR2 U2608 (.A(n2666),
	.B(n2078),
	.OUT(n1880));
   XOR2 U2609 (.A(n2670),
	.B(n2079),
	.OUT(n1878));
   XOR2 U2610 (.A(n2674),
	.B(n2080),
	.OUT(n1876));
   XOR2 U2611 (.A(n2678),
	.B(n2081),
	.OUT(n1874));
   XOR2 U2612 (.A(n2682),
	.B(n2082),
	.OUT(n1872));
   XOR2 U2613 (.A(n2686),
	.B(n2083),
	.OUT(n1870));
   XOR2 U2614 (.A(n2690),
	.B(n2084),
	.OUT(n1868));
   XOR2 U2615 (.A(n2694),
	.B(n2085),
	.OUT(n1866));
   XOR2 U2616 (.A(n2698),
	.B(n2086),
	.OUT(n1864));
   XOR2 U2617 (.A(n2815),
	.B(n2702),
	.OUT(n218));
   inverter U2618 (.IN(n741),
	.OUT(n1743));
   inverter U2619 (.IN(n738),
	.OUT(n2709));
   XOR2 U2620 (.A(n2708),
	.B(n2089),
	.OUT(n1914));
   XOR2 U2621 (.A(n2711),
	.B(n2090),
	.OUT(n1912));
   XOR2 U2622 (.A(n2715),
	.B(n2091),
	.OUT(n1910));
   XOR2 U2623 (.A(n2719),
	.B(n2092),
	.OUT(n1908));
   XOR2 U2624 (.A(n2723),
	.B(n2093),
	.OUT(n1906));
   XOR2 U2625 (.A(n2727),
	.B(n2094),
	.OUT(n1904));
   XOR2 U2626 (.A(n2731),
	.B(n2095),
	.OUT(n1902));
   XOR2 U2627 (.A(n2735),
	.B(n2096),
	.OUT(n1900));
   XOR2 U2628 (.A(n2739),
	.B(n2097),
	.OUT(n1898));
   XOR2 U2629 (.A(n2743),
	.B(n2098),
	.OUT(n1896));
   XOR2 U2630 (.A(n2747),
	.B(n2099),
	.OUT(n1894));
   XOR2 U2631 (.A(n2751),
	.B(n2100),
	.OUT(n1892));
   XOR2 U2632 (.A(n2816),
	.B(n2755),
	.OUT(n228));
   XOR2 U2633 (.A(n748),
	.B(\mult_21_3/ab[2][3] ),
	.OUT(n245));
   XOR2 U2634 (.A(n752),
	.B(\mult_21_3/ab[2][4] ),
	.OUT(n242));
   XOR2 U2635 (.A(n2138),
	.B(n771),
	.OUT(n236));
   XOR2 U2636 (.A(\mult_21_3/ab[2][7] ),
	.B(n781),
	.OUT(n2760));
   XOR2 U2637 (.A(\mult_21_3/ab[3][7] ),
	.B(n793),
	.OUT(n2817));
   XOR2 U2638 (.A(n744),
	.B(\mult_21_3/ab[2][2] ),
	.OUT(n262));
   XOR2 U2639 (.A(n802),
	.B(\mult_21_3/ab[2][1] ),
	.OUT(n271));
   XOR2 U2640 (.A(\mult_21_3/ab[4][7] ),
	.B(\mult_21_3/ab[5][6] ),
	.OUT(n2763));
   XOR2 U2641 (.A(\mult_21_3/ab[5][7] ),
	.B(n835),
	.OUT(n2764));
   XOR2 U2642 (.A(\mult_21_3/ab[6][7] ),
	.B(\mult_21_3/ab[7][6] ),
	.OUT(n2765));
   XOR2 U2643 (.A(n848),
	.B(\mult_21_2/ab[2][3] ),
	.OUT(n300));
   XOR2 U2644 (.A(n852),
	.B(\mult_21_2/ab[2][4] ),
	.OUT(n297));
   XOR2 U2645 (.A(n2133),
	.B(n871),
	.OUT(n291));
   XOR2 U2646 (.A(\mult_21_2/ab[2][7] ),
	.B(n881),
	.OUT(n2766));
   XOR2 U2647 (.A(\mult_21_2/ab[3][7] ),
	.B(n893),
	.OUT(n2818));
   XOR2 U2648 (.A(n844),
	.B(\mult_21_2/ab[2][2] ),
	.OUT(n317));
   XOR2 U2649 (.A(n902),
	.B(\mult_21_2/ab[2][1] ),
	.OUT(n326));
   XOR2 U2650 (.A(\mult_21_2/ab[4][7] ),
	.B(\mult_21_2/ab[5][6] ),
	.OUT(n2769));
   XOR2 U2651 (.A(\mult_21_2/ab[5][7] ),
	.B(n935),
	.OUT(n2770));
   XOR2 U2652 (.A(\mult_21_2/ab[6][7] ),
	.B(\mult_21_2/ab[7][6] ),
	.OUT(n2771));
   XOR2 U2653 (.A(n948),
	.B(\mult_21/ab[2][3] ),
	.OUT(n355));
   XOR2 U2654 (.A(n952),
	.B(\mult_21/ab[2][4] ),
	.OUT(n352));
   XOR2 U2655 (.A(n2129),
	.B(n971),
	.OUT(n346));
   XOR2 U2656 (.A(\mult_21/ab[2][7] ),
	.B(n981),
	.OUT(n2772));
   XOR2 U2657 (.A(\mult_21/ab[3][7] ),
	.B(n993),
	.OUT(n2819));
   XOR2 U2658 (.A(n944),
	.B(\mult_21/ab[2][2] ),
	.OUT(n372));
   XOR2 U2659 (.A(n1002),
	.B(\mult_21/ab[2][1] ),
	.OUT(n381));
   XOR2 U2660 (.A(\mult_21/ab[4][7] ),
	.B(\mult_21/ab[5][6] ),
	.OUT(n2775));
   XOR2 U2661 (.A(\mult_21/ab[5][7] ),
	.B(n1035),
	.OUT(n2776));
   XOR2 U2662 (.A(\mult_21/ab[6][7] ),
	.B(\mult_21/ab[7][6] ),
	.OUT(n2777));
   XOR2 U2663 (.A(n1048),
	.B(\mult_20_3/ab[2][3] ),
	.OUT(n410));
   XOR2 U2664 (.A(n1052),
	.B(\mult_20_3/ab[2][4] ),
	.OUT(n407));
   XOR2 U2665 (.A(n2125),
	.B(n1071),
	.OUT(n401));
   XOR2 U2666 (.A(\mult_20_3/ab[2][7] ),
	.B(n1081),
	.OUT(n2778));
   XOR2 U2667 (.A(\mult_20_3/ab[3][7] ),
	.B(n1093),
	.OUT(n2820));
   XOR2 U2668 (.A(n1044),
	.B(\mult_20_3/ab[2][2] ),
	.OUT(n427));
   XOR2 U2669 (.A(n1102),
	.B(\mult_20_3/ab[2][1] ),
	.OUT(n436));
   XOR2 U2670 (.A(\mult_20_3/ab[4][7] ),
	.B(\mult_20_3/ab[5][6] ),
	.OUT(n2781));
   XOR2 U2671 (.A(\mult_20_3/ab[5][7] ),
	.B(n1135),
	.OUT(n2782));
   XOR2 U2672 (.A(\mult_20_3/ab[6][7] ),
	.B(\mult_20_3/ab[7][6] ),
	.OUT(n2783));
   XOR2 U2673 (.A(n1148),
	.B(\mult_20_2/ab[2][3] ),
	.OUT(n465));
   XOR2 U2674 (.A(n1152),
	.B(\mult_20_2/ab[2][4] ),
	.OUT(n462));
   XOR2 U2675 (.A(n2120),
	.B(n1171),
	.OUT(n456));
   XOR2 U2676 (.A(\mult_20_2/ab[2][7] ),
	.B(n1181),
	.OUT(n2784));
   XOR2 U2677 (.A(\mult_20_2/ab[3][7] ),
	.B(n1193),
	.OUT(n2821));
   XOR2 U2678 (.A(n1144),
	.B(\mult_20_2/ab[2][2] ),
	.OUT(n482));
   XOR2 U2679 (.A(n1202),
	.B(\mult_20_2/ab[2][1] ),
	.OUT(n491));
   XOR2 U2680 (.A(\mult_20_2/ab[4][7] ),
	.B(\mult_20_2/ab[5][6] ),
	.OUT(n2787));
   XOR2 U2681 (.A(\mult_20_2/ab[5][7] ),
	.B(n1235),
	.OUT(n2788));
   XOR2 U2682 (.A(\mult_20_2/ab[6][7] ),
	.B(\mult_20_2/ab[7][6] ),
	.OUT(n2789));
   XOR2 U2683 (.A(n1248),
	.B(\mult_20/ab[2][3] ),
	.OUT(n520));
   XOR2 U2684 (.A(n1252),
	.B(\mult_20/ab[2][4] ),
	.OUT(n517));
   XOR2 U2685 (.A(n2116),
	.B(n1271),
	.OUT(n511));
   XOR2 U2686 (.A(\mult_20/ab[2][7] ),
	.B(n1281),
	.OUT(n2790));
   XOR2 U2687 (.A(\mult_20/ab[3][7] ),
	.B(n1293),
	.OUT(n2822));
   XOR2 U2688 (.A(n1244),
	.B(\mult_20/ab[2][2] ),
	.OUT(n537));
   XOR2 U2689 (.A(n1302),
	.B(\mult_20/ab[2][1] ),
	.OUT(n546));
   XOR2 U2690 (.A(\mult_20/ab[4][7] ),
	.B(\mult_20/ab[5][6] ),
	.OUT(n2793));
   XOR2 U2691 (.A(\mult_20/ab[5][7] ),
	.B(n1335),
	.OUT(n2794));
   XOR2 U2692 (.A(\mult_20/ab[6][7] ),
	.B(\mult_20/ab[7][6] ),
	.OUT(n2795));
   XOR2 U2693 (.A(n1348),
	.B(\mult_19_3/ab[2][3] ),
	.OUT(n575));
   XOR2 U2694 (.A(n1352),
	.B(\mult_19_3/ab[2][4] ),
	.OUT(n572));
   XOR2 U2695 (.A(n2112),
	.B(n1371),
	.OUT(n566));
   XOR2 U2696 (.A(\mult_19_3/ab[2][7] ),
	.B(n1381),
	.OUT(n2796));
   XOR2 U2697 (.A(\mult_19_3/ab[3][7] ),
	.B(n1393),
	.OUT(n2823));
   XOR2 U2698 (.A(n1344),
	.B(\mult_19_3/ab[2][2] ),
	.OUT(n592));
   XOR2 U2699 (.A(n1402),
	.B(\mult_19_3/ab[2][1] ),
	.OUT(n601));
   XOR2 U2700 (.A(\mult_19_3/ab[4][7] ),
	.B(\mult_19_3/ab[5][6] ),
	.OUT(n2799));
   XOR2 U2701 (.A(\mult_19_3/ab[5][7] ),
	.B(n1435),
	.OUT(n2800));
   XOR2 U2702 (.A(\mult_19_3/ab[6][7] ),
	.B(\mult_19_3/ab[7][6] ),
	.OUT(n2801));
   XOR2 U2703 (.A(n1448),
	.B(\mult_19_2/ab[2][3] ),
	.OUT(n630));
   XOR2 U2704 (.A(n1452),
	.B(\mult_19_2/ab[2][4] ),
	.OUT(n627));
   XOR2 U2705 (.A(n2107),
	.B(n1471),
	.OUT(n621));
   XOR2 U2706 (.A(\mult_19_2/ab[2][7] ),
	.B(n1481),
	.OUT(n2802));
   XOR2 U2707 (.A(\mult_19_2/ab[3][7] ),
	.B(n1493),
	.OUT(n2824));
   XOR2 U2708 (.A(n1444),
	.B(\mult_19_2/ab[2][2] ),
	.OUT(n647));
   XOR2 U2709 (.A(n1502),
	.B(\mult_19_2/ab[2][1] ),
	.OUT(n656));
   XOR2 U2710 (.A(\mult_19_2/ab[4][7] ),
	.B(\mult_19_2/ab[5][6] ),
	.OUT(n2805));
   XOR2 U2711 (.A(\mult_19_2/ab[5][7] ),
	.B(n1535),
	.OUT(n2806));
   XOR2 U2712 (.A(\mult_19_2/ab[6][7] ),
	.B(\mult_19_2/ab[7][6] ),
	.OUT(n2807));
   XOR2 U2713 (.A(n1548),
	.B(\mult_19/ab[2][3] ),
	.OUT(n685));
   XOR2 U2714 (.A(n1552),
	.B(\mult_19/ab[2][4] ),
	.OUT(n682));
   XOR2 U2715 (.A(n2103),
	.B(n1571),
	.OUT(n676));
   XOR2 U2716 (.A(\mult_19/ab[2][7] ),
	.B(n1581),
	.OUT(n2808));
   XOR2 U2717 (.A(\mult_19/ab[3][7] ),
	.B(n1593),
	.OUT(n2825));
   XOR2 U2718 (.A(n1544),
	.B(\mult_19/ab[2][2] ),
	.OUT(n702));
   XOR2 U2719 (.A(n1602),
	.B(\mult_19/ab[2][1] ),
	.OUT(n711));
   XOR2 U2720 (.A(\mult_19/ab[4][7] ),
	.B(\mult_19/ab[5][6] ),
	.OUT(n2811));
   XOR2 U2721 (.A(\mult_19/ab[5][7] ),
	.B(n1635),
	.OUT(n2812));
   XOR2 U2722 (.A(\mult_19/ab[6][7] ),
	.B(\mult_19/ab[7][6] ),
	.OUT(n2813));
   XOR2 U2723 (.A(n2111),
	.B(n726),
	.OUT(n731));
   XOR2 U2724 (.A(N31),
	.B(N15),
	.OUT(n2814));
   XOR2 U2725 (.A(n2137),
	.B(n732),
	.OUT(n737));
   XOR2 U2726 (.A(N191),
	.B(N175),
	.OUT(n2815));
   XOR2 U2727 (.A(n2124),
	.B(n738),
	.OUT(n743));
   XOR2 U2728 (.A(N111),
	.B(N95),
	.OUT(n2816));
   inverter U2729 (.IN(n2142),
	.OUT(n2144));
   inverter U2730 (.IN(n2151),
	.OUT(n792));
   inverter U2731 (.IN(n2147),
	.OUT(n796));
   inverter U2732 (.IN(n788),
	.OUT(n2149));
   inverter U2733 (.IN(n2165),
	.OUT(n2166));
   inverter U2734 (.IN(n2184),
	.OUT(n2185));
   inverter U2735 (.IN(n190),
	.OUT(\mult_21_3/A2[11] ));
   inverter U2736 (.IN(n2190),
	.OUT(n2192));
   inverter U2737 (.IN(n2193),
	.OUT(n2195));
   inverter U2738 (.IN(n2202),
	.OUT(n892));
   inverter U2739 (.IN(n2198),
	.OUT(n896));
   inverter U2740 (.IN(n888),
	.OUT(n2200));
   inverter U2741 (.IN(n2216),
	.OUT(n2217));
   inverter U2742 (.IN(n2235),
	.OUT(n2236));
   inverter U2743 (.IN(n175),
	.OUT(\mult_21_2/A2[11] ));
   inverter U2744 (.IN(n2241),
	.OUT(n2243));
   inverter U2745 (.IN(n2244),
	.OUT(n2246));
   inverter U2746 (.IN(n2253),
	.OUT(n992));
   inverter U2747 (.IN(n2249),
	.OUT(n996));
   inverter U2748 (.IN(n988),
	.OUT(n2251));
   inverter U2749 (.IN(n2267),
	.OUT(n2268));
   inverter U2750 (.IN(n2286),
	.OUT(n2287));
   inverter U2751 (.IN(n160),
	.OUT(\mult_21/A2[11] ));
   inverter U2752 (.IN(n2292),
	.OUT(n2294));
   inverter U2753 (.IN(n2295),
	.OUT(n2297));
   inverter U2754 (.IN(n2304),
	.OUT(n1092));
   inverter U2755 (.IN(n2300),
	.OUT(n1096));
   inverter U2756 (.IN(n1088),
	.OUT(n2302));
   inverter U2757 (.IN(n2318),
	.OUT(n2319));
   inverter U2758 (.IN(n2337),
	.OUT(n2338));
   inverter U2759 (.IN(n145),
	.OUT(\mult_20_3/A2[11] ));
   inverter U2760 (.IN(n2343),
	.OUT(n2345));
   inverter U2761 (.IN(n2346),
	.OUT(n2348));
   inverter U2762 (.IN(n2355),
	.OUT(n1192));
   inverter U2763 (.IN(n2351),
	.OUT(n1196));
   inverter U2764 (.IN(n1188),
	.OUT(n2353));
   inverter U2765 (.IN(n2369),
	.OUT(n2370));
   inverter U2766 (.IN(n2388),
	.OUT(n2389));
   inverter U2767 (.IN(n130),
	.OUT(\mult_20_2/A2[11] ));
   inverter U2768 (.IN(n2394),
	.OUT(n2396));
   inverter U2769 (.IN(n2397),
	.OUT(n2399));
   inverter U2770 (.IN(n2406),
	.OUT(n1292));
   inverter U2771 (.IN(n2402),
	.OUT(n1296));
   inverter U2772 (.IN(n1288),
	.OUT(n2404));
   inverter U2773 (.IN(n2420),
	.OUT(n2421));
   inverter U2774 (.IN(n2439),
	.OUT(n2440));
   inverter U2775 (.IN(n115),
	.OUT(\mult_20/A2[11] ));
   inverter U2776 (.IN(n2445),
	.OUT(n2447));
   inverter U2777 (.IN(n2448),
	.OUT(n2450));
   inverter U2778 (.IN(n2457),
	.OUT(n1392));
   inverter U2779 (.IN(n2453),
	.OUT(n1396));
   inverter U2780 (.IN(n1388),
	.OUT(n2455));
   inverter U2781 (.IN(n2471),
	.OUT(n2472));
   inverter U2782 (.IN(n2490),
	.OUT(n2491));
   inverter U2783 (.IN(n100),
	.OUT(\mult_19_3/A2[11] ));
   inverter U2784 (.IN(n2496),
	.OUT(n2498));
   inverter U2785 (.IN(n2499),
	.OUT(n2501));
   inverter U2786 (.IN(n2508),
	.OUT(n1492));
   inverter U2787 (.IN(n2504),
	.OUT(n1496));
   inverter U2788 (.IN(n1488),
	.OUT(n2506));
   inverter U2789 (.IN(n2522),
	.OUT(n2523));
   inverter U2790 (.IN(n2541),
	.OUT(n2542));
   inverter U2791 (.IN(n85),
	.OUT(\mult_19_2/A2[11] ));
   inverter U2792 (.IN(n2547),
	.OUT(n2549));
   inverter U2793 (.IN(n2550),
	.OUT(n2552));
   inverter U2794 (.IN(n2559),
	.OUT(n1592));
   inverter U2795 (.IN(n2555),
	.OUT(n1596));
   inverter U2796 (.IN(n1588),
	.OUT(n2557));
   inverter U2797 (.IN(n2573),
	.OUT(n2574));
   inverter U2798 (.IN(n2592),
	.OUT(n2593));
   inverter U2799 (.IN(n70),
	.OUT(\mult_19/A2[11] ));
   inverter U2800 (.IN(n2598),
	.OUT(n2600));
   inverter U2801 (.IN(n2604),
	.OUT(n2606));
   inverter U2802 (.IN(n2651),
	.OUT(n1650));
   inverter U2803 (.IN(n2657),
	.OUT(n2659));
   inverter U2804 (.IN(n2704),
	.OUT(n1698));
   inverter U2805 (.IN(n2710),
	.OUT(n2712));
   inverter U2806 (.IN(n2757),
	.OUT(n1746));
   inverter U2807 (.IN(n2155),
	.OUT(n758));
   inverter U2808 (.IN(n2156),
	.OUT(n768));
   inverter U2809 (.IN(\mult_21_3/ab[4][3] ),
	.OUT(n777));
   inverter U2810 (.IN(n2157),
	.OUT(n780));
   inverter U2811 (.IN(\mult_21_3/ab[3][5] ),
	.OUT(n785));
   inverter U2812 (.IN(n2159),
	.OUT(n2160));
   inverter U2813 (.IN(\mult_21_3/ab[6][3] ),
	.OUT(n800));
   inverter U2814 (.IN(n2167),
	.OUT(n820));
   inverter U2815 (.IN(n2168),
	.OUT(n823));
   inverter U2816 (.IN(n2169),
	.OUT(n825));
   inverter U2817 (.IN(n2170),
	.OUT(n828));
   inverter U2818 (.IN(n2171),
	.OUT(n830));
   inverter U2819 (.IN(\mult_21_3/ab[7][4] ),
	.OUT(n2189));
   inverter U2820 (.IN(n2206),
	.OUT(n858));
   inverter U2821 (.IN(n2207),
	.OUT(n868));
   inverter U2822 (.IN(\mult_21_2/ab[4][3] ),
	.OUT(n877));
   inverter U2823 (.IN(n2208),
	.OUT(n880));
   inverter U2824 (.IN(\mult_21_2/ab[3][5] ),
	.OUT(n885));
   inverter U2825 (.IN(n2210),
	.OUT(n2211));
   inverter U2826 (.IN(\mult_21_2/ab[6][3] ),
	.OUT(n900));
   inverter U2827 (.IN(n2218),
	.OUT(n920));
   inverter U2828 (.IN(n2219),
	.OUT(n923));
   inverter U2829 (.IN(n2220),
	.OUT(n925));
   inverter U2830 (.IN(n2221),
	.OUT(n928));
   inverter U2831 (.IN(n2222),
	.OUT(n930));
   inverter U2832 (.IN(\mult_21_2/ab[7][4] ),
	.OUT(n2240));
   inverter U2833 (.IN(n2257),
	.OUT(n958));
   inverter U2834 (.IN(n2258),
	.OUT(n968));
   inverter U2835 (.IN(\mult_21/ab[4][3] ),
	.OUT(n977));
   inverter U2836 (.IN(n2259),
	.OUT(n980));
   inverter U2837 (.IN(\mult_21/ab[3][5] ),
	.OUT(n985));
   inverter U2838 (.IN(n2261),
	.OUT(n2262));
   inverter U2839 (.IN(\mult_21/ab[6][3] ),
	.OUT(n1000));
   inverter U2840 (.IN(n2269),
	.OUT(n1020));
   inverter U2841 (.IN(n2270),
	.OUT(n1023));
   inverter U2842 (.IN(n2271),
	.OUT(n1025));
   inverter U2843 (.IN(n2272),
	.OUT(n1028));
   inverter U2844 (.IN(n2273),
	.OUT(n1030));
   inverter U2845 (.IN(\mult_21/ab[7][4] ),
	.OUT(n2291));
   inverter U2846 (.IN(n2308),
	.OUT(n1058));
   inverter U2847 (.IN(n2309),
	.OUT(n1068));
   inverter U2848 (.IN(\mult_20_3/ab[4][3] ),
	.OUT(n1077));
   inverter U2849 (.IN(n2310),
	.OUT(n1080));
   inverter U2850 (.IN(\mult_20_3/ab[3][5] ),
	.OUT(n1085));
   inverter U2851 (.IN(n2312),
	.OUT(n2313));
   inverter U2852 (.IN(\mult_20_3/ab[6][3] ),
	.OUT(n1100));
   inverter U2853 (.IN(n2320),
	.OUT(n1120));
   inverter U2854 (.IN(n2321),
	.OUT(n1123));
   inverter U2855 (.IN(n2322),
	.OUT(n1125));
   inverter U2856 (.IN(n2323),
	.OUT(n1128));
   inverter U2857 (.IN(n2324),
	.OUT(n1130));
   inverter U2858 (.IN(\mult_20_3/ab[7][4] ),
	.OUT(n2342));
   inverter U2859 (.IN(n2359),
	.OUT(n1158));
   inverter U2860 (.IN(n2360),
	.OUT(n1168));
   inverter U2861 (.IN(\mult_20_2/ab[4][3] ),
	.OUT(n1177));
   inverter U2862 (.IN(n2361),
	.OUT(n1180));
   inverter U2863 (.IN(\mult_20_2/ab[3][5] ),
	.OUT(n1185));
   inverter U2864 (.IN(n2363),
	.OUT(n2364));
   inverter U2865 (.IN(\mult_20_2/ab[6][3] ),
	.OUT(n1200));
   inverter U2866 (.IN(n2371),
	.OUT(n1220));
   inverter U2867 (.IN(n2372),
	.OUT(n1223));
   inverter U2868 (.IN(n2373),
	.OUT(n1225));
   inverter U2869 (.IN(n2374),
	.OUT(n1228));
   inverter U2870 (.IN(n2375),
	.OUT(n1230));
   inverter U2871 (.IN(\mult_20_2/ab[7][4] ),
	.OUT(n2393));
   inverter U2872 (.IN(n2410),
	.OUT(n1258));
   inverter U2873 (.IN(n2411),
	.OUT(n1268));
   inverter U2874 (.IN(\mult_20/ab[4][3] ),
	.OUT(n1277));
   inverter U2875 (.IN(n2412),
	.OUT(n1280));
   inverter U2876 (.IN(\mult_20/ab[3][5] ),
	.OUT(n1285));
   inverter U2877 (.IN(n2414),
	.OUT(n2415));
   inverter U2878 (.IN(\mult_20/ab[6][3] ),
	.OUT(n1300));
   inverter U2879 (.IN(n2422),
	.OUT(n1320));
   inverter U2880 (.IN(n2423),
	.OUT(n1323));
   inverter U2881 (.IN(n2424),
	.OUT(n1325));
   inverter U2882 (.IN(n2425),
	.OUT(n1328));
   inverter U2883 (.IN(n2426),
	.OUT(n1330));
   inverter U2884 (.IN(\mult_20/ab[7][4] ),
	.OUT(n2444));
   inverter U2885 (.IN(n2461),
	.OUT(n1358));
   inverter U2886 (.IN(n2462),
	.OUT(n1368));
   inverter U2887 (.IN(\mult_19_3/ab[4][3] ),
	.OUT(n1377));
   inverter U2888 (.IN(n2463),
	.OUT(n1380));
   inverter U2889 (.IN(\mult_19_3/ab[3][5] ),
	.OUT(n1385));
   inverter U2890 (.IN(n2465),
	.OUT(n2466));
   inverter U2891 (.IN(\mult_19_3/ab[6][3] ),
	.OUT(n1400));
   inverter U2892 (.IN(n2473),
	.OUT(n1420));
   inverter U2893 (.IN(n2474),
	.OUT(n1423));
   inverter U2894 (.IN(n2475),
	.OUT(n1425));
   inverter U2895 (.IN(n2476),
	.OUT(n1428));
   inverter U2896 (.IN(n2477),
	.OUT(n1430));
   inverter U2897 (.IN(\mult_19_3/ab[7][4] ),
	.OUT(n2495));
   inverter U2898 (.IN(n2512),
	.OUT(n1458));
   inverter U2899 (.IN(n2513),
	.OUT(n1468));
   inverter U2900 (.IN(\mult_19_2/ab[4][3] ),
	.OUT(n1477));
   inverter U2901 (.IN(n2514),
	.OUT(n1480));
   inverter U2902 (.IN(\mult_19_2/ab[3][5] ),
	.OUT(n1485));
   inverter U2903 (.IN(n2516),
	.OUT(n2517));
   inverter U2904 (.IN(\mult_19_2/ab[6][3] ),
	.OUT(n1500));
   inverter U2905 (.IN(n2524),
	.OUT(n1520));
   inverter U2906 (.IN(n2525),
	.OUT(n1523));
   inverter U2907 (.IN(n2526),
	.OUT(n1525));
   inverter U2908 (.IN(n2527),
	.OUT(n1528));
   inverter U2909 (.IN(n2528),
	.OUT(n1530));
   inverter U2910 (.IN(\mult_19_2/ab[7][4] ),
	.OUT(n2546));
   inverter U2911 (.IN(n2563),
	.OUT(n1558));
   inverter U2912 (.IN(n2564),
	.OUT(n1568));
   inverter U2913 (.IN(\mult_19/ab[4][3] ),
	.OUT(n1577));
   inverter U2914 (.IN(n2565),
	.OUT(n1580));
   inverter U2915 (.IN(\mult_19/ab[3][5] ),
	.OUT(n1585));
   inverter U2916 (.IN(n2567),
	.OUT(n2568));
   inverter U2917 (.IN(\mult_19/ab[6][3] ),
	.OUT(n1600));
   inverter U2918 (.IN(n2575),
	.OUT(n1620));
   inverter U2919 (.IN(n2576),
	.OUT(n1623));
   inverter U2920 (.IN(n2577),
	.OUT(n1625));
   inverter U2921 (.IN(n2578),
	.OUT(n1628));
   inverter U2922 (.IN(n2579),
	.OUT(n1630));
   inverter U2923 (.IN(\mult_19/ab[7][4] ),
	.OUT(n2597));
   inverter U2924 (.IN(n2153),
	.OUT(n747));
   inverter U2925 (.IN(n2154),
	.OUT(n751));
   inverter U2926 (.IN(n2152),
	.OUT(n801));
   inverter U2927 (.IN(\mult_21_3/ab[4][1] ),
	.OUT(n810));
   inverter U2928 (.IN(n2183),
	.OUT(n841));
   inverter U2929 (.IN(n2186),
	.OUT(n843));
   inverter U2930 (.IN(n2204),
	.OUT(n847));
   inverter U2931 (.IN(n2205),
	.OUT(n851));
   inverter U2932 (.IN(n2203),
	.OUT(n901));
   inverter U2933 (.IN(\mult_21_2/ab[4][1] ),
	.OUT(n910));
   inverter U2934 (.IN(n2234),
	.OUT(n941));
   inverter U2935 (.IN(n2237),
	.OUT(n943));
   inverter U2936 (.IN(n2255),
	.OUT(n947));
   inverter U2937 (.IN(n2256),
	.OUT(n951));
   inverter U2938 (.IN(n2254),
	.OUT(n1001));
   inverter U2939 (.IN(\mult_21/ab[4][1] ),
	.OUT(n1010));
   inverter U2940 (.IN(n2285),
	.OUT(n1041));
   inverter U2941 (.IN(n2288),
	.OUT(n1043));
   inverter U2942 (.IN(n2306),
	.OUT(n1047));
   inverter U2943 (.IN(n2307),
	.OUT(n1051));
   inverter U2944 (.IN(n2305),
	.OUT(n1101));
   inverter U2945 (.IN(\mult_20_3/ab[4][1] ),
	.OUT(n1110));
   inverter U2946 (.IN(n2336),
	.OUT(n1141));
   inverter U2947 (.IN(n2339),
	.OUT(n1143));
   inverter U2948 (.IN(n2357),
	.OUT(n1147));
   inverter U2949 (.IN(n2358),
	.OUT(n1151));
   inverter U2950 (.IN(n2356),
	.OUT(n1201));
   inverter U2951 (.IN(\mult_20_2/ab[4][1] ),
	.OUT(n1210));
   inverter U2952 (.IN(n2387),
	.OUT(n1241));
   inverter U2953 (.IN(n2390),
	.OUT(n1243));
   inverter U2954 (.IN(n2408),
	.OUT(n1247));
   inverter U2955 (.IN(n2409),
	.OUT(n1251));
   inverter U2956 (.IN(n2407),
	.OUT(n1301));
   inverter U2957 (.IN(\mult_20/ab[4][1] ),
	.OUT(n1310));
   inverter U2958 (.IN(n2438),
	.OUT(n1341));
   inverter U2959 (.IN(n2441),
	.OUT(n1343));
   inverter U2960 (.IN(n2459),
	.OUT(n1347));
   inverter U2961 (.IN(n2460),
	.OUT(n1351));
   inverter U2962 (.IN(n2458),
	.OUT(n1401));
   inverter U2963 (.IN(\mult_19_3/ab[4][1] ),
	.OUT(n1410));
   inverter U2964 (.IN(n2489),
	.OUT(n1441));
   inverter U2965 (.IN(n2492),
	.OUT(n1443));
   inverter U2966 (.IN(n2510),
	.OUT(n1447));
   inverter U2967 (.IN(n2511),
	.OUT(n1451));
   inverter U2968 (.IN(n2509),
	.OUT(n1501));
   inverter U2969 (.IN(\mult_19_2/ab[4][1] ),
	.OUT(n1510));
   inverter U2970 (.IN(n2540),
	.OUT(n1541));
   inverter U2971 (.IN(n2543),
	.OUT(n1543));
   inverter U2972 (.IN(n2561),
	.OUT(n1547));
   inverter U2973 (.IN(n2562),
	.OUT(n1551));
   inverter U2974 (.IN(n2560),
	.OUT(n1601));
   inverter U2975 (.IN(\mult_19/ab[4][1] ),
	.OUT(n1610));
   inverter U2976 (.IN(n2591),
	.OUT(n1641));
   inverter U2977 (.IN(n2594),
	.OUT(n1643));
   inverter U2978 (.IN(n1662),
	.OUT(n1667));
   inverter U2979 (.IN(n1670),
	.OUT(n1675));
   inverter U2980 (.IN(n1678),
	.OUT(n1683));
   inverter U2981 (.IN(n1710),
	.OUT(n1715));
   inverter U2982 (.IN(n1718),
	.OUT(n1723));
   inverter U2983 (.IN(n1726),
	.OUT(n1731));
   inverter U2984 (.IN(n1758),
	.OUT(n1763));
   inverter U2985 (.IN(n1766),
	.OUT(n1771));
   inverter U2986 (.IN(n1774),
	.OUT(n1779));
   inverter U2987 (.IN(n803),
	.OUT(n2161));
   inverter U2988 (.IN(n2163),
	.OUT(n813));
   inverter U2989 (.IN(n903),
	.OUT(n2212));
   inverter U2990 (.IN(n2214),
	.OUT(n913));
   inverter U2991 (.IN(n1003),
	.OUT(n2263));
   inverter U2992 (.IN(n2265),
	.OUT(n1013));
   inverter U2993 (.IN(n1103),
	.OUT(n2314));
   inverter U2994 (.IN(n2316),
	.OUT(n1113));
   inverter U2995 (.IN(n1203),
	.OUT(n2365));
   inverter U2996 (.IN(n2367),
	.OUT(n1213));
   inverter U2997 (.IN(n1303),
	.OUT(n2416));
   inverter U2998 (.IN(n2418),
	.OUT(n1313));
   inverter U2999 (.IN(n1403),
	.OUT(n2467));
   inverter U3000 (.IN(n2469),
	.OUT(n1413));
   inverter U3001 (.IN(n1503),
	.OUT(n2518));
   inverter U3002 (.IN(n2520),
	.OUT(n1513));
   inverter U3003 (.IN(n1603),
	.OUT(n2569));
   inverter U3004 (.IN(n2571),
	.OUT(n1613));
   inverter U3005 (.IN(n1652),
	.OUT(n2653));
   inverter U3006 (.IN(n1700),
	.OUT(n2706));
   inverter U3007 (.IN(n1748),
	.OUT(n2759));
   inverter U3008 (.IN(n754),
	.OUT(n2150));
   inverter U3009 (.IN(\mult_21_3/ab[2][5] ),
	.OUT(n771));
   inverter U3010 (.IN(n761),
	.OUT(n2148));
   inverter U3011 (.IN(\mult_21_3/ab[2][1] ),
	.OUT(n804));
   inverter U3012 (.IN(\mult_21_3/ab[5][5] ),
	.OUT(n1924));
   inverter U3013 (.IN(n854),
	.OUT(n2201));
   inverter U3014 (.IN(\mult_21_2/ab[2][5] ),
	.OUT(n871));
   inverter U3015 (.IN(n861),
	.OUT(n2199));
   inverter U3016 (.IN(\mult_21_2/ab[2][1] ),
	.OUT(n904));
   inverter U3017 (.IN(\mult_21_2/ab[5][5] ),
	.OUT(n1940));
   inverter U3018 (.IN(n954),
	.OUT(n2252));
   inverter U3019 (.IN(\mult_21/ab[2][5] ),
	.OUT(n971));
   inverter U3020 (.IN(n961),
	.OUT(n2250));
   inverter U3021 (.IN(\mult_21/ab[2][1] ),
	.OUT(n1004));
   inverter U3022 (.IN(\mult_21/ab[5][5] ),
	.OUT(n1956));
   inverter U3023 (.IN(n1054),
	.OUT(n2303));
   inverter U3024 (.IN(\mult_20_3/ab[2][5] ),
	.OUT(n1071));
   inverter U3025 (.IN(n1061),
	.OUT(n2301));
   inverter U3026 (.IN(\mult_20_3/ab[2][1] ),
	.OUT(n1104));
   inverter U3027 (.IN(\mult_20_3/ab[5][5] ),
	.OUT(n1972));
   inverter U3028 (.IN(n1154),
	.OUT(n2354));
   inverter U3029 (.IN(\mult_20_2/ab[2][5] ),
	.OUT(n1171));
   inverter U3030 (.IN(n1161),
	.OUT(n2352));
   inverter U3031 (.IN(\mult_20_2/ab[2][1] ),
	.OUT(n1204));
   inverter U3032 (.IN(\mult_20_2/ab[5][5] ),
	.OUT(n1988));
   inverter U3033 (.IN(n1254),
	.OUT(n2405));
   inverter U3034 (.IN(\mult_20/ab[2][5] ),
	.OUT(n1271));
   inverter U3035 (.IN(n1261),
	.OUT(n2403));
   inverter U3036 (.IN(\mult_20/ab[2][1] ),
	.OUT(n1304));
   inverter U3037 (.IN(\mult_20/ab[5][5] ),
	.OUT(n2004));
   inverter U3038 (.IN(n1354),
	.OUT(n2456));
   inverter U3039 (.IN(\mult_19_3/ab[2][5] ),
	.OUT(n1371));
   inverter U3040 (.IN(n1361),
	.OUT(n2454));
   inverter U3041 (.IN(\mult_19_3/ab[2][1] ),
	.OUT(n1404));
   inverter U3042 (.IN(\mult_19_3/ab[5][5] ),
	.OUT(n2020));
   inverter U3043 (.IN(n1454),
	.OUT(n2507));
   inverter U3044 (.IN(\mult_19_2/ab[2][5] ),
	.OUT(n1471));
   inverter U3045 (.IN(n1461),
	.OUT(n2505));
   inverter U3046 (.IN(\mult_19_2/ab[2][1] ),
	.OUT(n1504));
   inverter U3047 (.IN(\mult_19_2/ab[5][5] ),
	.OUT(n2036));
   inverter U3048 (.IN(n1554),
	.OUT(n2558));
   inverter U3049 (.IN(\mult_19/ab[2][5] ),
	.OUT(n1571));
   inverter U3050 (.IN(n1561),
	.OUT(n2556));
   inverter U3051 (.IN(\mult_19/ab[2][1] ),
	.OUT(n1604));
   inverter U3052 (.IN(\mult_19/ab[5][5] ),
	.OUT(n2052));
   inverter U3053 (.IN(n1655),
	.OUT(n1659));
   inverter U3054 (.IN(n1666),
	.OUT(n1671));
   inverter U3055 (.IN(n1674),
	.OUT(n1679));
   inverter U3056 (.IN(n1682),
	.OUT(n1687));
   inverter U3057 (.IN(n1703),
	.OUT(n1707));
   inverter U3058 (.IN(n1714),
	.OUT(n1719));
   inverter U3059 (.IN(n1722),
	.OUT(n1727));
   inverter U3060 (.IN(n1730),
	.OUT(n1735));
   inverter U3061 (.IN(n1751),
	.OUT(n1755));
   inverter U3062 (.IN(n1762),
	.OUT(n1767));
   inverter U3063 (.IN(n1770),
	.OUT(n1775));
   inverter U3064 (.IN(n1778),
	.OUT(n1783));
   inverter U3065 (.IN(\mult_21_3/ab[2][3] ),
	.OUT(n755));
   inverter U3066 (.IN(\mult_21_3/ab[2][4] ),
	.OUT(n762));
   inverter U3067 (.IN(n774),
	.OUT(n789));
   inverter U3068 (.IN(n2817),
	.OUT(n2761));
   inverter U3069 (.IN(n2191),
	.OUT(n258));
   inverter U3070 (.IN(n2762),
	.OUT(n200));
   inverter U3071 (.IN(n2179),
	.OUT(n2181));
   inverter U3072 (.IN(n2180),
	.OUT(n2182));
   inverter U3073 (.IN(\mult_21_2/ab[2][3] ),
	.OUT(n855));
   inverter U3074 (.IN(\mult_21_2/ab[2][4] ),
	.OUT(n862));
   inverter U3075 (.IN(n874),
	.OUT(n889));
   inverter U3076 (.IN(n2818),
	.OUT(n2767));
   inverter U3077 (.IN(n2242),
	.OUT(n313));
   inverter U3078 (.IN(n2768),
	.OUT(n185));
   inverter U3079 (.IN(n2230),
	.OUT(n2232));
   inverter U3080 (.IN(n2231),
	.OUT(n2233));
   inverter U3081 (.IN(\mult_21/ab[2][3] ),
	.OUT(n955));
   inverter U3082 (.IN(\mult_21/ab[2][4] ),
	.OUT(n962));
   inverter U3083 (.IN(n974),
	.OUT(n989));
   inverter U3084 (.IN(n2819),
	.OUT(n2773));
   inverter U3085 (.IN(n2293),
	.OUT(n368));
   inverter U3086 (.IN(n2774),
	.OUT(n170));
   inverter U3087 (.IN(n2281),
	.OUT(n2283));
   inverter U3088 (.IN(n2282),
	.OUT(n2284));
   inverter U3089 (.IN(\mult_20_3/ab[2][3] ),
	.OUT(n1055));
   inverter U3090 (.IN(\mult_20_3/ab[2][4] ),
	.OUT(n1062));
   inverter U3091 (.IN(n1074),
	.OUT(n1089));
   inverter U3092 (.IN(n2820),
	.OUT(n2779));
   inverter U3093 (.IN(n2344),
	.OUT(n423));
   inverter U3094 (.IN(n2780),
	.OUT(n155));
   inverter U3095 (.IN(n2332),
	.OUT(n2334));
   inverter U3096 (.IN(n2333),
	.OUT(n2335));
   inverter U3097 (.IN(\mult_20_2/ab[2][3] ),
	.OUT(n1155));
   inverter U3098 (.IN(\mult_20_2/ab[2][4] ),
	.OUT(n1162));
   inverter U3099 (.IN(n1174),
	.OUT(n1189));
   inverter U3100 (.IN(n2821),
	.OUT(n2785));
   inverter U3101 (.IN(n2395),
	.OUT(n478));
   inverter U3102 (.IN(n2786),
	.OUT(n140));
   inverter U3103 (.IN(n2383),
	.OUT(n2385));
   inverter U3104 (.IN(n2384),
	.OUT(n2386));
   inverter U3105 (.IN(\mult_20/ab[2][3] ),
	.OUT(n1255));
   inverter U3106 (.IN(\mult_20/ab[2][4] ),
	.OUT(n1262));
   inverter U3107 (.IN(n1274),
	.OUT(n1289));
   inverter U3108 (.IN(n2822),
	.OUT(n2791));
   inverter U3109 (.IN(n2446),
	.OUT(n533));
   inverter U3110 (.IN(n2792),
	.OUT(n125));
   inverter U3111 (.IN(n2434),
	.OUT(n2436));
   inverter U3112 (.IN(n2435),
	.OUT(n2437));
   inverter U3113 (.IN(\mult_19_3/ab[2][3] ),
	.OUT(n1355));
   inverter U3114 (.IN(\mult_19_3/ab[2][4] ),
	.OUT(n1362));
   inverter U3115 (.IN(n1374),
	.OUT(n1389));
   inverter U3116 (.IN(n2823),
	.OUT(n2797));
   inverter U3117 (.IN(n2497),
	.OUT(n588));
   inverter U3118 (.IN(n2798),
	.OUT(n110));
   inverter U3119 (.IN(n2485),
	.OUT(n2487));
   inverter U3120 (.IN(n2486),
	.OUT(n2488));
   inverter U3121 (.IN(\mult_19_2/ab[2][3] ),
	.OUT(n1455));
   inverter U3122 (.IN(\mult_19_2/ab[2][4] ),
	.OUT(n1462));
   inverter U3123 (.IN(n1474),
	.OUT(n1489));
   inverter U3124 (.IN(n2824),
	.OUT(n2803));
   inverter U3125 (.IN(n2548),
	.OUT(n643));
   inverter U3126 (.IN(n2804),
	.OUT(n95));
   inverter U3127 (.IN(n2536),
	.OUT(n2538));
   inverter U3128 (.IN(n2537),
	.OUT(n2539));
   inverter U3129 (.IN(\mult_19/ab[2][3] ),
	.OUT(n1555));
   inverter U3130 (.IN(\mult_19/ab[2][4] ),
	.OUT(n1562));
   inverter U3131 (.IN(n1574),
	.OUT(n1589));
   inverter U3132 (.IN(n2825),
	.OUT(n2809));
   inverter U3133 (.IN(n2599),
	.OUT(n698));
   inverter U3134 (.IN(n2810),
	.OUT(n80));
   inverter U3135 (.IN(n2587),
	.OUT(n2589));
   inverter U3136 (.IN(n2588),
	.OUT(n2590));
   inverter U3137 (.IN(n2605),
	.OUT(n2608));
   inverter U3138 (.IN(n2607),
	.OUT(n2610));
   inverter U3139 (.IN(n2609),
	.OUT(n2612));
   inverter U3140 (.IN(n2611),
	.OUT(n2614));
   inverter U3141 (.IN(n2613),
	.OUT(n2616));
   inverter U3142 (.IN(n2615),
	.OUT(n2618));
   inverter U3143 (.IN(n2617),
	.OUT(n2620));
   inverter U3144 (.IN(n2619),
	.OUT(n2622));
   inverter U3145 (.IN(n2621),
	.OUT(n2624));
   inverter U3146 (.IN(n2623),
	.OUT(n2626));
   inverter U3147 (.IN(n2625),
	.OUT(n2628));
   inverter U3148 (.IN(n2627),
	.OUT(n2630));
   inverter U3149 (.IN(n2629),
	.OUT(n2632));
   inverter U3150 (.IN(n2631),
	.OUT(n2634));
   inverter U3151 (.IN(n2633),
	.OUT(n2636));
   inverter U3152 (.IN(n2635),
	.OUT(n2638));
   inverter U3153 (.IN(n2637),
	.OUT(n2640));
   inverter U3154 (.IN(n2639),
	.OUT(n2642));
   inverter U3155 (.IN(n2641),
	.OUT(n2644));
   inverter U3156 (.IN(n2643),
	.OUT(n2646));
   inverter U3157 (.IN(n2645),
	.OUT(n2648));
   inverter U3158 (.IN(n2647),
	.OUT(n2650));
   inverter U3159 (.IN(n2649),
	.OUT(n202));
   inverter U3160 (.IN(n201),
	.OUT(n204));
   inverter U3161 (.IN(n2652),
	.OUT(n1653));
   inverter U3162 (.IN(n1658),
	.OUT(n1663));
   inverter U3163 (.IN(n1686),
	.OUT(n1690));
   inverter U3164 (.IN(n2658),
	.OUT(n2661));
   inverter U3165 (.IN(n2660),
	.OUT(n2663));
   inverter U3166 (.IN(n2662),
	.OUT(n2665));
   inverter U3167 (.IN(n2664),
	.OUT(n2667));
   inverter U3168 (.IN(n2666),
	.OUT(n2669));
   inverter U3169 (.IN(n2668),
	.OUT(n2671));
   inverter U3170 (.IN(n2670),
	.OUT(n2673));
   inverter U3171 (.IN(n2672),
	.OUT(n2675));
   inverter U3172 (.IN(n2674),
	.OUT(n2677));
   inverter U3173 (.IN(n2676),
	.OUT(n2679));
   inverter U3174 (.IN(n2678),
	.OUT(n2681));
   inverter U3175 (.IN(n2680),
	.OUT(n2683));
   inverter U3176 (.IN(n2682),
	.OUT(n2685));
   inverter U3177 (.IN(n2684),
	.OUT(n2687));
   inverter U3178 (.IN(n2686),
	.OUT(n2689));
   inverter U3179 (.IN(n2688),
	.OUT(n2691));
   inverter U3180 (.IN(n2690),
	.OUT(n2693));
   inverter U3181 (.IN(n2692),
	.OUT(n2695));
   inverter U3182 (.IN(n2694),
	.OUT(n2697));
   inverter U3183 (.IN(n2696),
	.OUT(n2699));
   inverter U3184 (.IN(n2698),
	.OUT(n2701));
   inverter U3185 (.IN(n2700),
	.OUT(n2703));
   inverter U3186 (.IN(n2702),
	.OUT(n212));
   inverter U3187 (.IN(n211),
	.OUT(n214));
   inverter U3188 (.IN(n2705),
	.OUT(n1701));
   inverter U3189 (.IN(n1706),
	.OUT(n1711));
   inverter U3190 (.IN(n1734),
	.OUT(n1738));
   inverter U3191 (.IN(n2711),
	.OUT(n2714));
   inverter U3192 (.IN(n2713),
	.OUT(n2716));
   inverter U3193 (.IN(n2715),
	.OUT(n2718));
   inverter U3194 (.IN(n2717),
	.OUT(n2720));
   inverter U3195 (.IN(n2719),
	.OUT(n2722));
   inverter U3196 (.IN(n2721),
	.OUT(n2724));
   inverter U3197 (.IN(n2723),
	.OUT(n2726));
   inverter U3198 (.IN(n2725),
	.OUT(n2728));
   inverter U3199 (.IN(n2727),
	.OUT(n2730));
   inverter U3200 (.IN(n2729),
	.OUT(n2732));
   inverter U3201 (.IN(n2731),
	.OUT(n2734));
   inverter U3202 (.IN(n2733),
	.OUT(n2736));
   inverter U3203 (.IN(n2735),
	.OUT(n2738));
   inverter U3204 (.IN(n2737),
	.OUT(n2740));
   inverter U3205 (.IN(n2739),
	.OUT(n2742));
   inverter U3206 (.IN(n2741),
	.OUT(n2744));
   inverter U3207 (.IN(n2743),
	.OUT(n2746));
   inverter U3208 (.IN(n2745),
	.OUT(n2748));
   inverter U3209 (.IN(n2747),
	.OUT(n2750));
   inverter U3210 (.IN(n2749),
	.OUT(n2752));
   inverter U3211 (.IN(n2751),
	.OUT(n2754));
   inverter U3212 (.IN(n2753),
	.OUT(n2756));
   inverter U3213 (.IN(n2755),
	.OUT(n222));
   inverter U3214 (.IN(n221),
	.OUT(n224));
   inverter U3215 (.IN(n2758),
	.OUT(n1749));
   inverter U3216 (.IN(n1754),
	.OUT(n1759));
   inverter U3217 (.IN(n1782),
	.OUT(n1786));
   inverter U3218 (.IN(\mult_19/A1[0] ),
	.OUT(n2826));
   inverter U3219 (.IN(n2827),
	.OUT(N3));
   inverter U3220 (.IN(\mult_19/A1[1] ),
	.OUT(n2828));
   inverter U3221 (.IN(n2829),
	.OUT(N4));
   inverter U3222 (.IN(\mult_19/A1[2] ),
	.OUT(n2830));
   inverter U3223 (.IN(n2831),
	.OUT(N5));
   inverter U3224 (.IN(\mult_19/A1[3] ),
	.OUT(n2832));
   inverter U3225 (.IN(n2833),
	.OUT(N6));
   inverter U3226 (.IN(\mult_19/A1[4] ),
	.OUT(n2834));
   inverter U3227 (.IN(n2835),
	.OUT(N7));
   inverter U3228 (.IN(\mult_19/A1[5] ),
	.OUT(n2836));
   inverter U3229 (.IN(n2837),
	.OUT(N8));
   inverter U3230 (.IN(\mult_19/A1[6] ),
	.OUT(n2838));
   inverter U3231 (.IN(n2839),
	.OUT(N9));
   inverter U3232 (.IN(\mult_19/A1[7] ),
	.OUT(n2840));
   inverter U3233 (.IN(\mult_19/A2[7] ),
	.OUT(n2841));
   inverter U3234 (.IN(n2842),
	.OUT(N10));
   inverter U3235 (.IN(\mult_19/A1[8] ),
	.OUT(n2843));
   inverter U3236 (.IN(\mult_19/A2[8] ),
	.OUT(n2844));
   inverter U3237 (.IN(n2845),
	.OUT(\mult_19/FS_1/PG_int[0][2][0] ));
   inverter U3238 (.IN(\mult_19/A1[9] ),
	.OUT(n2846));
   inverter U3239 (.IN(\mult_19/A2[9] ),
	.OUT(n2847));
   inverter U3240 (.IN(n2848),
	.OUT(\mult_19/FS_1/PG_int[0][2][1] ));
   inverter U3241 (.IN(n2849),
	.OUT(\mult_19/FS_1/TEMP_P[0][2][1] ));
   inverter U3242 (.IN(\mult_19/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2850));
   inverter U3243 (.IN(\mult_19/A1[10] ),
	.OUT(n2851));
   inverter U3244 (.IN(\mult_19/A2[10] ),
	.OUT(n2852));
   inverter U3245 (.IN(n2853),
	.OUT(\mult_19/FS_1/PG_int[0][2][2] ));
   inverter U3246 (.IN(n2854),
	.OUT(\mult_19/FS_1/TEMP_P[0][2][2] ));
   inverter U3247 (.IN(\mult_19/FS_1/TEMP_G[0][2][1] ),
	.OUT(n2855));
   inverter U3248 (.IN(\mult_19/FS_1/C[1][2][1] ),
	.OUT(n2856));
   inverter U3249 (.IN(\mult_19/FS_1/P[0][2][1] ),
	.OUT(n2857));
   inverter U3250 (.IN(\mult_19/A1[11] ),
	.OUT(n2858));
   inverter U3251 (.IN(\mult_19/A2[11] ),
	.OUT(n2859));
   inverter U3252 (.IN(n2860),
	.OUT(\mult_19/FS_1/PG_int[0][2][3] ));
   inverter U3253 (.IN(\mult_19/FS_1/TEMP_G[0][2][2] ),
	.OUT(n2861));
   inverter U3254 (.IN(\mult_19/FS_1/P[0][2][3] ),
	.OUT(n2862));
   inverter U3255 (.IN(\mult_19/FS_1/C[1][2][2] ),
	.OUT(n2863));
   inverter U3256 (.IN(\mult_19/FS_1/P[0][2][2] ),
	.OUT(n2864));
   inverter U3257 (.IN(\mult_19/A1[12] ),
	.OUT(n2865));
   inverter U3258 (.IN(\mult_19/A2[12] ),
	.OUT(n2866));
   inverter U3259 (.IN(n2867),
	.OUT(\mult_19/FS_1/PG_int[0][3][0] ));
   inverter U3260 (.IN(\mult_19/A2[13] ),
	.OUT(n2868));
   inverter U3261 (.IN(n2869),
	.OUT(\mult_19/FS_1/PG_int[0][3][1] ));
   inverter U3262 (.IN(\mult_19/FS_1/C[1][3][0] ),
	.OUT(n2870));
   inverter U3263 (.IN(\mult_19/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2871));
   inverter U3264 (.IN(\mult_19/FS_1/G[1][0][1] ),
	.OUT(n2872));
   inverter U3265 (.IN(\mult_19/FS_1/C[1][2][0] ),
	.OUT(n2873));
   inverter U3266 (.IN(\mult_19/FS_1/G[1][0][2] ),
	.OUT(n2875));
   inverter U3267 (.IN(\mult_19_2/A1[0] ),
	.OUT(n2876));
   inverter U3268 (.IN(n2877),
	.OUT(N19));
   inverter U3269 (.IN(\mult_19_2/A1[1] ),
	.OUT(n2878));
   inverter U3270 (.IN(n2879),
	.OUT(N20));
   inverter U3271 (.IN(\mult_19_2/A1[2] ),
	.OUT(n2880));
   inverter U3272 (.IN(n2881),
	.OUT(N21));
   inverter U3273 (.IN(\mult_19_2/A1[3] ),
	.OUT(n2882));
   inverter U3274 (.IN(n2883),
	.OUT(N22));
   inverter U3275 (.IN(\mult_19_2/A1[4] ),
	.OUT(n2884));
   inverter U3276 (.IN(n2885),
	.OUT(N23));
   inverter U3277 (.IN(\mult_19_2/A1[5] ),
	.OUT(n2886));
   inverter U3278 (.IN(n2887),
	.OUT(N24));
   inverter U3279 (.IN(\mult_19_2/A1[6] ),
	.OUT(n2888));
   inverter U3280 (.IN(n2889),
	.OUT(N25));
   inverter U3281 (.IN(\mult_19_2/A1[7] ),
	.OUT(n2890));
   inverter U3282 (.IN(\mult_19_2/A2[7] ),
	.OUT(n2891));
   inverter U3283 (.IN(n2892),
	.OUT(N26));
   inverter U3284 (.IN(\mult_19_2/A1[8] ),
	.OUT(n2893));
   inverter U3285 (.IN(\mult_19_2/A2[8] ),
	.OUT(n2894));
   inverter U3286 (.IN(n2895),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][0] ));
   inverter U3287 (.IN(\mult_19_2/A1[9] ),
	.OUT(n2896));
   inverter U3288 (.IN(\mult_19_2/A2[9] ),
	.OUT(n2897));
   inverter U3289 (.IN(n2898),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][1] ));
   inverter U3290 (.IN(n2899),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][2][1] ));
   inverter U3291 (.IN(\mult_19_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2900));
   inverter U3292 (.IN(\mult_19_2/A1[10] ),
	.OUT(n2901));
   inverter U3293 (.IN(\mult_19_2/A2[10] ),
	.OUT(n2902));
   inverter U3294 (.IN(n2903),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][2] ));
   inverter U3295 (.IN(n2904),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][2][2] ));
   inverter U3296 (.IN(\mult_19_2/FS_1/TEMP_G[0][2][1] ),
	.OUT(n2905));
   inverter U3297 (.IN(\mult_19_2/FS_1/C[1][2][1] ),
	.OUT(n2906));
   inverter U3298 (.IN(\mult_19_2/FS_1/P[0][2][1] ),
	.OUT(n2907));
   inverter U3299 (.IN(\mult_19_2/A1[11] ),
	.OUT(n2908));
   inverter U3300 (.IN(\mult_19_2/A2[11] ),
	.OUT(n2909));
   inverter U3301 (.IN(n2910),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][3] ));
   inverter U3302 (.IN(\mult_19_2/FS_1/TEMP_G[0][2][2] ),
	.OUT(n2911));
   inverter U3303 (.IN(\mult_19_2/FS_1/P[0][2][3] ),
	.OUT(n2912));
   inverter U3304 (.IN(\mult_19_2/FS_1/C[1][2][2] ),
	.OUT(n2913));
   inverter U3305 (.IN(\mult_19_2/FS_1/P[0][2][2] ),
	.OUT(n2914));
   inverter U3306 (.IN(\mult_19_2/A1[12] ),
	.OUT(n2915));
   inverter U3307 (.IN(\mult_19_2/A2[12] ),
	.OUT(n2916));
   inverter U3308 (.IN(n2917),
	.OUT(\mult_19_2/FS_1/PG_int[0][3][0] ));
   inverter U3309 (.IN(\mult_19_2/A2[13] ),
	.OUT(n2918));
   inverter U3310 (.IN(n2919),
	.OUT(\mult_19_2/FS_1/PG_int[0][3][1] ));
   inverter U3311 (.IN(\mult_19_2/FS_1/C[1][3][0] ),
	.OUT(n2920));
   inverter U3312 (.IN(\mult_19_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2921));
   inverter U3313 (.IN(\mult_19_2/FS_1/G[1][0][1] ),
	.OUT(n2922));
   inverter U3314 (.IN(\mult_19_2/FS_1/C[1][2][0] ),
	.OUT(n2923));
   inverter U3315 (.IN(\mult_19_2/FS_1/G[1][0][2] ),
	.OUT(n2925));
   inverter U3316 (.IN(\mult_19_3/A1[0] ),
	.OUT(n2926));
   inverter U3317 (.IN(n2927),
	.OUT(N51));
   inverter U3318 (.IN(\mult_19_3/A1[1] ),
	.OUT(n2928));
   inverter U3319 (.IN(n2929),
	.OUT(N52));
   inverter U3320 (.IN(\mult_19_3/A1[2] ),
	.OUT(n2930));
   inverter U3321 (.IN(n2931),
	.OUT(N53));
   inverter U3322 (.IN(\mult_19_3/A1[3] ),
	.OUT(n2932));
   inverter U3323 (.IN(n2933),
	.OUT(N54));
   inverter U3324 (.IN(\mult_19_3/A1[4] ),
	.OUT(n2934));
   inverter U3325 (.IN(n2935),
	.OUT(N55));
   inverter U3326 (.IN(\mult_19_3/A1[5] ),
	.OUT(n2936));
   inverter U3327 (.IN(n2937),
	.OUT(N56));
   inverter U3328 (.IN(\mult_19_3/A1[6] ),
	.OUT(n2938));
   inverter U3329 (.IN(n2939),
	.OUT(N57));
   inverter U3330 (.IN(\mult_19_3/A1[7] ),
	.OUT(n2940));
   inverter U3331 (.IN(\mult_19_3/A2[7] ),
	.OUT(n2941));
   inverter U3332 (.IN(n2942),
	.OUT(N58));
   inverter U3333 (.IN(\mult_19_3/A1[8] ),
	.OUT(n2943));
   inverter U3334 (.IN(\mult_19_3/A2[8] ),
	.OUT(n2944));
   inverter U3335 (.IN(n2945),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][0] ));
   inverter U3336 (.IN(\mult_19_3/A1[9] ),
	.OUT(n2946));
   inverter U3337 (.IN(\mult_19_3/A2[9] ),
	.OUT(n2947));
   inverter U3338 (.IN(n2948),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][1] ));
   inverter U3339 (.IN(n2949),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][2][1] ));
   inverter U3340 (.IN(\mult_19_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2950));
   inverter U3341 (.IN(\mult_19_3/A1[10] ),
	.OUT(n2951));
   inverter U3342 (.IN(\mult_19_3/A2[10] ),
	.OUT(n2952));
   inverter U3343 (.IN(n2953),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][2] ));
   inverter U3344 (.IN(n2954),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][2][2] ));
   inverter U3345 (.IN(\mult_19_3/FS_1/TEMP_G[0][2][1] ),
	.OUT(n2955));
   inverter U3346 (.IN(\mult_19_3/FS_1/C[1][2][1] ),
	.OUT(n2956));
   inverter U3347 (.IN(\mult_19_3/FS_1/P[0][2][1] ),
	.OUT(n2957));
   inverter U3348 (.IN(\mult_19_3/A1[11] ),
	.OUT(n2958));
   inverter U3349 (.IN(\mult_19_3/A2[11] ),
	.OUT(n2959));
   inverter U3350 (.IN(n2960),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][3] ));
   inverter U3351 (.IN(\mult_19_3/FS_1/TEMP_G[0][2][2] ),
	.OUT(n2961));
   inverter U3352 (.IN(\mult_19_3/FS_1/P[0][2][3] ),
	.OUT(n2962));
   inverter U3353 (.IN(\mult_19_3/FS_1/C[1][2][2] ),
	.OUT(n2963));
   inverter U3354 (.IN(\mult_19_3/FS_1/P[0][2][2] ),
	.OUT(n2964));
   inverter U3355 (.IN(\mult_19_3/A1[12] ),
	.OUT(n2965));
   inverter U3356 (.IN(\mult_19_3/A2[12] ),
	.OUT(n2966));
   inverter U3357 (.IN(n2967),
	.OUT(\mult_19_3/FS_1/PG_int[0][3][0] ));
   inverter U3358 (.IN(\mult_19_3/A2[13] ),
	.OUT(n2968));
   inverter U3359 (.IN(n2969),
	.OUT(\mult_19_3/FS_1/PG_int[0][3][1] ));
   inverter U3360 (.IN(\mult_19_3/FS_1/C[1][3][0] ),
	.OUT(n2970));
   inverter U3361 (.IN(\mult_19_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2971));
   inverter U3362 (.IN(\mult_19_3/FS_1/G[1][0][1] ),
	.OUT(n2972));
   inverter U3363 (.IN(\mult_19_3/FS_1/C[1][2][0] ),
	.OUT(n2973));
   inverter U3364 (.IN(\mult_19_3/FS_1/G[1][0][2] ),
	.OUT(n2975));
   inverter U3365 (.IN(\mult_20/A1[0] ),
	.OUT(n2976));
   inverter U3366 (.IN(n2977),
	.OUT(N83));
   inverter U3367 (.IN(\mult_20/A1[1] ),
	.OUT(n2978));
   inverter U3368 (.IN(n2979),
	.OUT(N84));
   inverter U3369 (.IN(\mult_20/A1[2] ),
	.OUT(n2980));
   inverter U3370 (.IN(n2981),
	.OUT(N85));
   inverter U3371 (.IN(\mult_20/A1[3] ),
	.OUT(n2982));
   inverter U3372 (.IN(n2983),
	.OUT(N86));
   inverter U3373 (.IN(\mult_20/A1[4] ),
	.OUT(n2984));
   inverter U3374 (.IN(n2985),
	.OUT(N87));
   inverter U3375 (.IN(\mult_20/A1[5] ),
	.OUT(n2986));
   inverter U3376 (.IN(n2987),
	.OUT(N88));
   inverter U3377 (.IN(\mult_20/A1[6] ),
	.OUT(n2988));
   inverter U3378 (.IN(n2989),
	.OUT(N89));
   inverter U3379 (.IN(\mult_20/A1[7] ),
	.OUT(n2990));
   inverter U3380 (.IN(\mult_20/A2[7] ),
	.OUT(n2991));
   inverter U3381 (.IN(n2992),
	.OUT(N90));
   inverter U3382 (.IN(\mult_20/A1[8] ),
	.OUT(n2993));
   inverter U3383 (.IN(\mult_20/A2[8] ),
	.OUT(n2994));
   inverter U3384 (.IN(n2995),
	.OUT(\mult_20/FS_1/PG_int[0][2][0] ));
   inverter U3385 (.IN(\mult_20/A1[9] ),
	.OUT(n2996));
   inverter U3386 (.IN(\mult_20/A2[9] ),
	.OUT(n2997));
   inverter U3387 (.IN(n2998),
	.OUT(\mult_20/FS_1/PG_int[0][2][1] ));
   inverter U3388 (.IN(n2999),
	.OUT(\mult_20/FS_1/TEMP_P[0][2][1] ));
   inverter U3389 (.IN(\mult_20/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3000));
   inverter U3390 (.IN(\mult_20/A1[10] ),
	.OUT(n3001));
   inverter U3391 (.IN(\mult_20/A2[10] ),
	.OUT(n3002));
   inverter U3392 (.IN(n3003),
	.OUT(\mult_20/FS_1/PG_int[0][2][2] ));
   inverter U3393 (.IN(n3004),
	.OUT(\mult_20/FS_1/TEMP_P[0][2][2] ));
   inverter U3394 (.IN(\mult_20/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3005));
   inverter U3395 (.IN(\mult_20/FS_1/C[1][2][1] ),
	.OUT(n3006));
   inverter U3396 (.IN(\mult_20/FS_1/P[0][2][1] ),
	.OUT(n3007));
   inverter U3397 (.IN(\mult_20/A1[11] ),
	.OUT(n3008));
   inverter U3398 (.IN(\mult_20/A2[11] ),
	.OUT(n3009));
   inverter U3399 (.IN(n3010),
	.OUT(\mult_20/FS_1/PG_int[0][2][3] ));
   inverter U3400 (.IN(\mult_20/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3011));
   inverter U3401 (.IN(\mult_20/FS_1/P[0][2][3] ),
	.OUT(n3012));
   inverter U3402 (.IN(\mult_20/FS_1/C[1][2][2] ),
	.OUT(n3013));
   inverter U3403 (.IN(\mult_20/FS_1/P[0][2][2] ),
	.OUT(n3014));
   inverter U3404 (.IN(\mult_20/A1[12] ),
	.OUT(n3015));
   inverter U3405 (.IN(\mult_20/A2[12] ),
	.OUT(n3016));
   inverter U3406 (.IN(n3017),
	.OUT(\mult_20/FS_1/PG_int[0][3][0] ));
   inverter U3407 (.IN(\mult_20/A2[13] ),
	.OUT(n3018));
   inverter U3408 (.IN(n3019),
	.OUT(\mult_20/FS_1/PG_int[0][3][1] ));
   inverter U3409 (.IN(\mult_20/FS_1/C[1][3][0] ),
	.OUT(n3020));
   inverter U3410 (.IN(\mult_20/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3021));
   inverter U3411 (.IN(\mult_20/FS_1/G[1][0][1] ),
	.OUT(n3022));
   inverter U3412 (.IN(\mult_20/FS_1/C[1][2][0] ),
	.OUT(n3023));
   inverter U3413 (.IN(\mult_20/FS_1/G[1][0][2] ),
	.OUT(n3025));
   inverter U3414 (.IN(\mult_20_2/A1[0] ),
	.OUT(n3026));
   inverter U3415 (.IN(n3027),
	.OUT(N99));
   inverter U3416 (.IN(\mult_20_2/A1[1] ),
	.OUT(n3028));
   inverter U3417 (.IN(n3029),
	.OUT(N100));
   inverter U3418 (.IN(\mult_20_2/A1[2] ),
	.OUT(n3030));
   inverter U3419 (.IN(n3031),
	.OUT(N101));
   inverter U3420 (.IN(\mult_20_2/A1[3] ),
	.OUT(n3032));
   inverter U3421 (.IN(n3033),
	.OUT(N102));
   inverter U3422 (.IN(\mult_20_2/A1[4] ),
	.OUT(n3034));
   inverter U3423 (.IN(n3035),
	.OUT(N103));
   inverter U3424 (.IN(\mult_20_2/A1[5] ),
	.OUT(n3036));
   inverter U3425 (.IN(n3037),
	.OUT(N104));
   inverter U3426 (.IN(\mult_20_2/A1[6] ),
	.OUT(n3038));
   inverter U3427 (.IN(n3039),
	.OUT(N105));
   inverter U3428 (.IN(\mult_20_2/A1[7] ),
	.OUT(n3040));
   inverter U3429 (.IN(\mult_20_2/A2[7] ),
	.OUT(n3041));
   inverter U3430 (.IN(n3042),
	.OUT(N106));
   inverter U3431 (.IN(\mult_20_2/A1[8] ),
	.OUT(n3043));
   inverter U3432 (.IN(\mult_20_2/A2[8] ),
	.OUT(n3044));
   inverter U3433 (.IN(n3045),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][0] ));
   inverter U3434 (.IN(\mult_20_2/A1[9] ),
	.OUT(n3046));
   inverter U3435 (.IN(\mult_20_2/A2[9] ),
	.OUT(n3047));
   inverter U3436 (.IN(n3048),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][1] ));
   inverter U3437 (.IN(n3049),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][2][1] ));
   inverter U3438 (.IN(\mult_20_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3050));
   inverter U3439 (.IN(\mult_20_2/A1[10] ),
	.OUT(n3051));
   inverter U3440 (.IN(\mult_20_2/A2[10] ),
	.OUT(n3052));
   inverter U3441 (.IN(n3053),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][2] ));
   inverter U3442 (.IN(n3054),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][2][2] ));
   inverter U3443 (.IN(\mult_20_2/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3055));
   inverter U3444 (.IN(\mult_20_2/FS_1/C[1][2][1] ),
	.OUT(n3056));
   inverter U3445 (.IN(\mult_20_2/FS_1/P[0][2][1] ),
	.OUT(n3057));
   inverter U3446 (.IN(\mult_20_2/A1[11] ),
	.OUT(n3058));
   inverter U3447 (.IN(\mult_20_2/A2[11] ),
	.OUT(n3059));
   inverter U3448 (.IN(n3060),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][3] ));
   inverter U3449 (.IN(\mult_20_2/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3061));
   inverter U3450 (.IN(\mult_20_2/FS_1/P[0][2][3] ),
	.OUT(n3062));
   inverter U3451 (.IN(\mult_20_2/FS_1/C[1][2][2] ),
	.OUT(n3063));
   inverter U3452 (.IN(\mult_20_2/FS_1/P[0][2][2] ),
	.OUT(n3064));
   inverter U3453 (.IN(\mult_20_2/A1[12] ),
	.OUT(n3065));
   inverter U3454 (.IN(\mult_20_2/A2[12] ),
	.OUT(n3066));
   inverter U3455 (.IN(n3067),
	.OUT(\mult_20_2/FS_1/PG_int[0][3][0] ));
   inverter U3456 (.IN(\mult_20_2/A2[13] ),
	.OUT(n3068));
   inverter U3457 (.IN(n3069),
	.OUT(\mult_20_2/FS_1/PG_int[0][3][1] ));
   inverter U3458 (.IN(\mult_20_2/FS_1/C[1][3][0] ),
	.OUT(n3070));
   inverter U3459 (.IN(\mult_20_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3071));
   inverter U3460 (.IN(\mult_20_2/FS_1/G[1][0][1] ),
	.OUT(n3072));
   inverter U3461 (.IN(\mult_20_2/FS_1/C[1][2][0] ),
	.OUT(n3073));
   inverter U3462 (.IN(\mult_20_2/FS_1/G[1][0][2] ),
	.OUT(n3075));
   inverter U3463 (.IN(\mult_20_3/A1[0] ),
	.OUT(n3076));
   inverter U3464 (.IN(n3077),
	.OUT(N131));
   inverter U3465 (.IN(\mult_20_3/A1[1] ),
	.OUT(n3078));
   inverter U3466 (.IN(n3079),
	.OUT(N132));
   inverter U3467 (.IN(\mult_20_3/A1[2] ),
	.OUT(n3080));
   inverter U3468 (.IN(n3081),
	.OUT(N133));
   inverter U3469 (.IN(\mult_20_3/A1[3] ),
	.OUT(n3082));
   inverter U3470 (.IN(n3083),
	.OUT(N134));
   inverter U3471 (.IN(\mult_20_3/A1[4] ),
	.OUT(n3084));
   inverter U3472 (.IN(n3085),
	.OUT(N135));
   inverter U3473 (.IN(\mult_20_3/A1[5] ),
	.OUT(n3086));
   inverter U3474 (.IN(n3087),
	.OUT(N136));
   inverter U3475 (.IN(\mult_20_3/A1[6] ),
	.OUT(n3088));
   inverter U3476 (.IN(n3089),
	.OUT(N137));
   inverter U3477 (.IN(\mult_20_3/A1[7] ),
	.OUT(n3090));
   inverter U3478 (.IN(\mult_20_3/A2[7] ),
	.OUT(n3091));
   inverter U3479 (.IN(n3092),
	.OUT(N138));
   inverter U3480 (.IN(\mult_20_3/A1[8] ),
	.OUT(n3093));
   inverter U3481 (.IN(\mult_20_3/A2[8] ),
	.OUT(n3094));
   inverter U3482 (.IN(n3095),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][0] ));
   inverter U3483 (.IN(\mult_20_3/A1[9] ),
	.OUT(n3096));
   inverter U3484 (.IN(\mult_20_3/A2[9] ),
	.OUT(n3097));
   inverter U3485 (.IN(n3098),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][1] ));
   inverter U3486 (.IN(n3099),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][2][1] ));
   inverter U3487 (.IN(\mult_20_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3100));
   inverter U3488 (.IN(\mult_20_3/A1[10] ),
	.OUT(n3101));
   inverter U3489 (.IN(\mult_20_3/A2[10] ),
	.OUT(n3102));
   inverter U3490 (.IN(n3103),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][2] ));
   inverter U3491 (.IN(n3104),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][2][2] ));
   inverter U3492 (.IN(\mult_20_3/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3105));
   inverter U3493 (.IN(\mult_20_3/FS_1/C[1][2][1] ),
	.OUT(n3106));
   inverter U3494 (.IN(\mult_20_3/FS_1/P[0][2][1] ),
	.OUT(n3107));
   inverter U3495 (.IN(\mult_20_3/A1[11] ),
	.OUT(n3108));
   inverter U3496 (.IN(\mult_20_3/A2[11] ),
	.OUT(n3109));
   inverter U3497 (.IN(n3110),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][3] ));
   inverter U3498 (.IN(\mult_20_3/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3111));
   inverter U3499 (.IN(\mult_20_3/FS_1/P[0][2][3] ),
	.OUT(n3112));
   inverter U3500 (.IN(\mult_20_3/FS_1/C[1][2][2] ),
	.OUT(n3113));
   inverter U3501 (.IN(\mult_20_3/FS_1/P[0][2][2] ),
	.OUT(n3114));
   inverter U3502 (.IN(\mult_20_3/A1[12] ),
	.OUT(n3115));
   inverter U3503 (.IN(\mult_20_3/A2[12] ),
	.OUT(n3116));
   inverter U3504 (.IN(n3117),
	.OUT(\mult_20_3/FS_1/PG_int[0][3][0] ));
   inverter U3505 (.IN(\mult_20_3/A2[13] ),
	.OUT(n3118));
   inverter U3506 (.IN(n3119),
	.OUT(\mult_20_3/FS_1/PG_int[0][3][1] ));
   inverter U3507 (.IN(\mult_20_3/FS_1/C[1][3][0] ),
	.OUT(n3120));
   inverter U3508 (.IN(\mult_20_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3121));
   inverter U3509 (.IN(\mult_20_3/FS_1/G[1][0][1] ),
	.OUT(n3122));
   inverter U3510 (.IN(\mult_20_3/FS_1/C[1][2][0] ),
	.OUT(n3123));
   inverter U3511 (.IN(\mult_20_3/FS_1/G[1][0][2] ),
	.OUT(n3125));
   inverter U3512 (.IN(\mult_21/A1[0] ),
	.OUT(n3126));
   inverter U3513 (.IN(n3127),
	.OUT(N163));
   inverter U3514 (.IN(\mult_21/A1[1] ),
	.OUT(n3128));
   inverter U3515 (.IN(n3129),
	.OUT(N164));
   inverter U3516 (.IN(\mult_21/A1[2] ),
	.OUT(n3130));
   inverter U3517 (.IN(n3131),
	.OUT(N165));
   inverter U3518 (.IN(\mult_21/A1[3] ),
	.OUT(n3132));
   inverter U3519 (.IN(n3133),
	.OUT(N166));
   inverter U3520 (.IN(\mult_21/A1[4] ),
	.OUT(n3134));
   inverter U3521 (.IN(n3135),
	.OUT(N167));
   inverter U3522 (.IN(\mult_21/A1[5] ),
	.OUT(n3136));
   inverter U3523 (.IN(n3137),
	.OUT(N168));
   inverter U3524 (.IN(\mult_21/A1[6] ),
	.OUT(n3138));
   inverter U3525 (.IN(n3139),
	.OUT(N169));
   inverter U3526 (.IN(\mult_21/A1[7] ),
	.OUT(n3140));
   inverter U3527 (.IN(\mult_21/A2[7] ),
	.OUT(n3141));
   inverter U3528 (.IN(n3142),
	.OUT(N170));
   inverter U3529 (.IN(\mult_21/A1[8] ),
	.OUT(n3143));
   inverter U3530 (.IN(\mult_21/A2[8] ),
	.OUT(n3144));
   inverter U3531 (.IN(n3145),
	.OUT(\mult_21/FS_1/PG_int[0][2][0] ));
   inverter U3532 (.IN(\mult_21/A1[9] ),
	.OUT(n3146));
   inverter U3533 (.IN(\mult_21/A2[9] ),
	.OUT(n3147));
   inverter U3534 (.IN(n3148),
	.OUT(\mult_21/FS_1/PG_int[0][2][1] ));
   inverter U3535 (.IN(n3149),
	.OUT(\mult_21/FS_1/TEMP_P[0][2][1] ));
   inverter U3536 (.IN(\mult_21/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3150));
   inverter U3537 (.IN(\mult_21/A1[10] ),
	.OUT(n3151));
   inverter U3538 (.IN(\mult_21/A2[10] ),
	.OUT(n3152));
   inverter U3539 (.IN(n3153),
	.OUT(\mult_21/FS_1/PG_int[0][2][2] ));
   inverter U3540 (.IN(n3154),
	.OUT(\mult_21/FS_1/TEMP_P[0][2][2] ));
   inverter U3541 (.IN(\mult_21/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3155));
   inverter U3542 (.IN(\mult_21/FS_1/C[1][2][1] ),
	.OUT(n3156));
   inverter U3543 (.IN(\mult_21/FS_1/P[0][2][1] ),
	.OUT(n3157));
   inverter U3544 (.IN(\mult_21/A1[11] ),
	.OUT(n3158));
   inverter U3545 (.IN(\mult_21/A2[11] ),
	.OUT(n3159));
   inverter U3546 (.IN(n3160),
	.OUT(\mult_21/FS_1/PG_int[0][2][3] ));
   inverter U3547 (.IN(\mult_21/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3161));
   inverter U3548 (.IN(\mult_21/FS_1/P[0][2][3] ),
	.OUT(n3162));
   inverter U3549 (.IN(\mult_21/FS_1/C[1][2][2] ),
	.OUT(n3163));
   inverter U3550 (.IN(\mult_21/FS_1/P[0][2][2] ),
	.OUT(n3164));
   inverter U3551 (.IN(\mult_21/A1[12] ),
	.OUT(n3165));
   inverter U3552 (.IN(\mult_21/A2[12] ),
	.OUT(n3166));
   inverter U3553 (.IN(n3167),
	.OUT(\mult_21/FS_1/PG_int[0][3][0] ));
   inverter U3554 (.IN(\mult_21/A2[13] ),
	.OUT(n3168));
   inverter U3555 (.IN(n3169),
	.OUT(\mult_21/FS_1/PG_int[0][3][1] ));
   inverter U3556 (.IN(\mult_21/FS_1/C[1][3][0] ),
	.OUT(n3170));
   inverter U3557 (.IN(\mult_21/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3171));
   inverter U3558 (.IN(\mult_21/FS_1/G[1][0][1] ),
	.OUT(n3172));
   inverter U3559 (.IN(\mult_21/FS_1/C[1][2][0] ),
	.OUT(n3173));
   inverter U3560 (.IN(\mult_21/FS_1/G[1][0][2] ),
	.OUT(n3175));
   inverter U3561 (.IN(\mult_21_2/A1[0] ),
	.OUT(n3176));
   inverter U3562 (.IN(n3177),
	.OUT(N179));
   inverter U3563 (.IN(\mult_21_2/A1[1] ),
	.OUT(n3178));
   inverter U3564 (.IN(n3179),
	.OUT(N180));
   inverter U3565 (.IN(\mult_21_2/A1[2] ),
	.OUT(n3180));
   inverter U3566 (.IN(n3181),
	.OUT(N181));
   inverter U3567 (.IN(\mult_21_2/A1[3] ),
	.OUT(n3182));
   inverter U3568 (.IN(n3183),
	.OUT(N182));
   inverter U3569 (.IN(\mult_21_2/A1[4] ),
	.OUT(n3184));
   inverter U3570 (.IN(n3185),
	.OUT(N183));
   inverter U3571 (.IN(\mult_21_2/A1[5] ),
	.OUT(n3186));
   inverter U3572 (.IN(n3187),
	.OUT(N184));
   inverter U3573 (.IN(\mult_21_2/A1[6] ),
	.OUT(n3188));
   inverter U3574 (.IN(n3189),
	.OUT(N185));
   inverter U3575 (.IN(\mult_21_2/A1[7] ),
	.OUT(n3190));
   inverter U3576 (.IN(\mult_21_2/A2[7] ),
	.OUT(n3191));
   inverter U3577 (.IN(n3192),
	.OUT(N186));
   inverter U3578 (.IN(\mult_21_2/A1[8] ),
	.OUT(n3193));
   inverter U3579 (.IN(\mult_21_2/A2[8] ),
	.OUT(n3194));
   inverter U3580 (.IN(n3195),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][0] ));
   inverter U3581 (.IN(\mult_21_2/A1[9] ),
	.OUT(n3196));
   inverter U3582 (.IN(\mult_21_2/A2[9] ),
	.OUT(n3197));
   inverter U3583 (.IN(n3198),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][1] ));
   inverter U3584 (.IN(n3199),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][2][1] ));
   inverter U3585 (.IN(\mult_21_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3200));
   inverter U3586 (.IN(\mult_21_2/A1[10] ),
	.OUT(n3201));
   inverter U3587 (.IN(\mult_21_2/A2[10] ),
	.OUT(n3202));
   inverter U3588 (.IN(n3203),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][2] ));
   inverter U3589 (.IN(n3204),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][2][2] ));
   inverter U3590 (.IN(\mult_21_2/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3205));
   inverter U3591 (.IN(\mult_21_2/FS_1/C[1][2][1] ),
	.OUT(n3206));
   inverter U3592 (.IN(\mult_21_2/FS_1/P[0][2][1] ),
	.OUT(n3207));
   inverter U3593 (.IN(\mult_21_2/A1[11] ),
	.OUT(n3208));
   inverter U3594 (.IN(\mult_21_2/A2[11] ),
	.OUT(n3209));
   inverter U3595 (.IN(n3210),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][3] ));
   inverter U3596 (.IN(\mult_21_2/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3211));
   inverter U3597 (.IN(\mult_21_2/FS_1/P[0][2][3] ),
	.OUT(n3212));
   inverter U3598 (.IN(\mult_21_2/FS_1/C[1][2][2] ),
	.OUT(n3213));
   inverter U3599 (.IN(\mult_21_2/FS_1/P[0][2][2] ),
	.OUT(n3214));
   inverter U3600 (.IN(\mult_21_2/A1[12] ),
	.OUT(n3215));
   inverter U3601 (.IN(\mult_21_2/A2[12] ),
	.OUT(n3216));
   inverter U3602 (.IN(n3217),
	.OUT(\mult_21_2/FS_1/PG_int[0][3][0] ));
   inverter U3603 (.IN(\mult_21_2/A2[13] ),
	.OUT(n3218));
   inverter U3604 (.IN(n3219),
	.OUT(\mult_21_2/FS_1/PG_int[0][3][1] ));
   inverter U3605 (.IN(\mult_21_2/FS_1/C[1][3][0] ),
	.OUT(n3220));
   inverter U3606 (.IN(\mult_21_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3221));
   inverter U3607 (.IN(\mult_21_2/FS_1/G[1][0][1] ),
	.OUT(n3222));
   inverter U3608 (.IN(\mult_21_2/FS_1/C[1][2][0] ),
	.OUT(n3223));
   inverter U3609 (.IN(\mult_21_2/FS_1/G[1][0][2] ),
	.OUT(n3225));
   inverter U3610 (.IN(\mult_21_3/A1[0] ),
	.OUT(n3226));
   inverter U3611 (.IN(n3227),
	.OUT(N211));
   inverter U3612 (.IN(\mult_21_3/A1[1] ),
	.OUT(n3228));
   inverter U3613 (.IN(n3229),
	.OUT(N212));
   inverter U3614 (.IN(\mult_21_3/A1[2] ),
	.OUT(n3230));
   inverter U3615 (.IN(n3231),
	.OUT(N213));
   inverter U3616 (.IN(\mult_21_3/A1[3] ),
	.OUT(n3232));
   inverter U3617 (.IN(n3233),
	.OUT(N214));
   inverter U3618 (.IN(\mult_21_3/A1[4] ),
	.OUT(n3234));
   inverter U3619 (.IN(n3235),
	.OUT(N215));
   inverter U3620 (.IN(\mult_21_3/A1[5] ),
	.OUT(n3236));
   inverter U3621 (.IN(n3237),
	.OUT(N216));
   inverter U3622 (.IN(\mult_21_3/A1[6] ),
	.OUT(n3238));
   inverter U3623 (.IN(n3239),
	.OUT(N217));
   inverter U3624 (.IN(\mult_21_3/A1[7] ),
	.OUT(n3240));
   inverter U3625 (.IN(\mult_21_3/A2[7] ),
	.OUT(n3241));
   inverter U3626 (.IN(n3242),
	.OUT(N218));
   inverter U3627 (.IN(\mult_21_3/A1[8] ),
	.OUT(n3243));
   inverter U3628 (.IN(\mult_21_3/A2[8] ),
	.OUT(n3244));
   inverter U3629 (.IN(n3245),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][0] ));
   inverter U3630 (.IN(\mult_21_3/A1[9] ),
	.OUT(n3246));
   inverter U3631 (.IN(\mult_21_3/A2[9] ),
	.OUT(n3247));
   inverter U3632 (.IN(n3248),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][1] ));
   inverter U3633 (.IN(n3249),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][2][1] ));
   inverter U3634 (.IN(\mult_21_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3250));
   inverter U3635 (.IN(\mult_21_3/A1[10] ),
	.OUT(n3251));
   inverter U3636 (.IN(\mult_21_3/A2[10] ),
	.OUT(n3252));
   inverter U3637 (.IN(n3253),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][2] ));
   inverter U3638 (.IN(n3254),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][2][2] ));
   inverter U3639 (.IN(\mult_21_3/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3255));
   inverter U3640 (.IN(\mult_21_3/FS_1/C[1][2][1] ),
	.OUT(n3256));
   inverter U3641 (.IN(\mult_21_3/FS_1/P[0][2][1] ),
	.OUT(n3257));
   inverter U3642 (.IN(\mult_21_3/A1[11] ),
	.OUT(n3258));
   inverter U3643 (.IN(\mult_21_3/A2[11] ),
	.OUT(n3259));
   inverter U3644 (.IN(n3260),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][3] ));
   inverter U3645 (.IN(\mult_21_3/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3261));
   inverter U3646 (.IN(\mult_21_3/FS_1/P[0][2][3] ),
	.OUT(n3262));
   inverter U3647 (.IN(\mult_21_3/FS_1/C[1][2][2] ),
	.OUT(n3263));
   inverter U3648 (.IN(\mult_21_3/FS_1/P[0][2][2] ),
	.OUT(n3264));
   inverter U3649 (.IN(\mult_21_3/A1[12] ),
	.OUT(n3265));
   inverter U3650 (.IN(\mult_21_3/A2[12] ),
	.OUT(n3266));
   inverter U3651 (.IN(n3267),
	.OUT(\mult_21_3/FS_1/PG_int[0][3][0] ));
   inverter U3652 (.IN(\mult_21_3/A2[13] ),
	.OUT(n3268));
   inverter U3653 (.IN(n3269),
	.OUT(\mult_21_3/FS_1/PG_int[0][3][1] ));
   inverter U3654 (.IN(\mult_21_3/FS_1/C[1][3][0] ),
	.OUT(n3270));
   inverter U3655 (.IN(\mult_21_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3271));
   inverter U3656 (.IN(\mult_21_3/FS_1/G[1][0][1] ),
	.OUT(n3272));
   inverter U3657 (.IN(\mult_21_3/FS_1/C[1][2][0] ),
	.OUT(n3273));
   inverter U3658 (.IN(\mult_21_3/FS_1/G[1][0][2] ),
	.OUT(n3275));
endmodule
