* File: Tri_INV.pex.sp
* Created: Tue Dec  3 01:49:17 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt Tri_INV  GND! OUT VDD! EN IN
* 
XD0_noxref GND! VDD! DIODENWX  AREA=7.4572e-12 PERIM=1.0942e-05
XMMN2 NET9 EN GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.924e-13 AS=1.17e-13
+ PD=1.78e-06 PS=9.7e-07 NRD=0.405769 NRS=0.407692 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.7e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=1.302e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.2338e-14 PANW9=0
+ PANW10=0
XMMN1 NET15 IN GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=9.334e-14 AS=1.17e-13
+ PD=8.79e-07 PS=9.7e-07 NRD=0.365385 NRS=0.457692 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=8.82e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=1.302e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.2338e-14 PANW9=0
+ PANW10=0
XMMN0 OUT EN NET15 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.9916e-13 AS=9.334e-14
+ PD=1.806e-06 PS=8.79e-07 NRD=0.425 NRS=0.325 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=1.303e-06 SB=3.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=1.302e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.2338e-14 PANW9=0 PANW10=0
XMMP2 NET9 EN VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.664e-13 AS=1.62e-13
+ PD=2.18e-06 PS=1.17e-06 NRD=0.280556 NRS=0.441667 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.7e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0
+ PANW3=3.038e-15 PANW4=3.1e-15 PANW5=3.1e-15 PANW6=4.364e-14 PANW7=1.96e-14
+ PANW8=1.24e-14 PANW9=4.402e-15 PANW10=3.605e-14
XMMP0 NET15 IN VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.2924e-13 AS=1.62e-13
+ PD=1.079e-06 PS=1.17e-06 NRD=0.261111 NRS=0.183333 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.82e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0
+ PANW3=3.038e-15 PANW4=3.1e-15 PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14
+ PANW8=1.24e-14 PANW9=4.9042e-14 PANW10=5.549e-14
XMMP1 OUT NET9 NET15 VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.7576e-13 AS=1.2924e-13
+ PD=2.206e-06 PS=1.079e-06 NRD=0.308333 NRS=0.2375 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.303e-06 SB=3.83e-07 SD=0 PANW1=0 PANW2=0
+ PANW3=3.038e-15 PANW4=3.1e-15 PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14
+ PANW8=1.24e-14 PANW9=4.9042e-14 PANW10=5.549e-14
*
.include "Tri_INV.pex.sp.TRI_INV.pxi"
*
.ends
*
*
