// Created by ihdl
module matrix_vector_mult (
	clk, 
	rst_n, 
	matrix00, 
	matrix01, 
	matrix02, 
	matrix10, 
	matrix11, 
	matrix12, 
	matrix20, 
	matrix21, 
	matrix22, 
	vector_0, 
	vector_1, 
	vector_2, 
	result_0, 
	result_1, 
	result_2);
   input clk;
   input rst_n;
   input [7:0] matrix00;
   input [7:0] matrix01;
   input [7:0] matrix02;
   input [7:0] matrix10;
   input [7:0] matrix11;
   input [7:0] matrix12;
   input [7:0] matrix20;
   input [7:0] matrix21;
   input [7:0] matrix22;
   input [7:0] vector_0;
   input [7:0] vector_1;
   input [7:0] vector_2;
   output [15:0] result_0;
   output [15:0] result_1;
   output [15:0] result_2;

   // Internal wires
   wire N0;
   wire N1;
   wire N3;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N49;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N67;
   wire N68;
   wire N69;
   wire N70;
   wire N71;
   wire N72;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N129;
   wire N131;
   wire N132;
   wire N133;
   wire N134;
   wire N135;
   wire N136;
   wire N137;
   wire N138;
   wire N139;
   wire N140;
   wire N141;
   wire N142;
   wire N143;
   wire N144;
   wire N145;
   wire N146;
   wire N147;
   wire N148;
   wire N149;
   wire N150;
   wire N151;
   wire N152;
   wire N153;
   wire N154;
   wire N155;
   wire N156;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N209;
   wire N211;
   wire N212;
   wire N213;
   wire N214;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N221;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N227;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N233;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N239;
   wire N240;
   wire n1;
   wire \mult_21_3/FS_1/C[1][2][0] ;
   wire \mult_21_3/FS_1/C[1][2][1] ;
   wire \mult_21_3/FS_1/C[1][2][2] ;
   wire \mult_21_3/FS_1/C[1][2][3] ;
   wire \mult_21_3/FS_1/C[1][3][0] ;
   wire \mult_21_3/FS_1/C[1][3][1] ;
   wire \mult_21_3/FS_1/P[0][0][1] ;
   wire \mult_21_3/FS_1/P[0][0][2] ;
   wire \mult_21_3/FS_1/P[0][0][3] ;
   wire \mult_21_3/FS_1/P[0][1][1] ;
   wire \mult_21_3/FS_1/P[0][1][2] ;
   wire \mult_21_3/FS_1/P[0][1][3] ;
   wire \mult_21_3/FS_1/P[0][2][1] ;
   wire \mult_21_3/FS_1/P[0][2][2] ;
   wire \mult_21_3/FS_1/P[0][2][3] ;
   wire \mult_21_3/FS_1/P[0][3][1] ;
   wire \mult_21_3/FS_1/TEMP_P[0][0][0] ;
   wire \mult_21_3/FS_1/TEMP_P[0][1][0] ;
   wire \mult_21_3/FS_1/TEMP_P[0][2][0] ;
   wire \mult_21_3/FS_1/TEMP_P[0][2][1] ;
   wire \mult_21_3/FS_1/TEMP_P[0][2][2] ;
   wire \mult_21_3/FS_1/TEMP_P[0][3][0] ;
   wire \mult_21_3/FS_1/G[1][0][1] ;
   wire \mult_21_3/FS_1/G[1][0][2] ;
   wire \mult_21_3/FS_1/TEMP_G[0][2][1] ;
   wire \mult_21_3/FS_1/TEMP_G[0][2][2] ;
   wire \mult_21_3/FS_1/G_n_int[0][1][3] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][0] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][1] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][2] ;
   wire \mult_21_3/FS_1/G_n_int[0][2][3] ;
   wire \mult_21_3/FS_1/G_n_int[0][3][0] ;
   wire \mult_21_3/FS_1/PG_int[0][2][0] ;
   wire \mult_21_3/FS_1/PG_int[0][2][1] ;
   wire \mult_21_3/FS_1/PG_int[0][2][2] ;
   wire \mult_21_3/FS_1/PG_int[0][2][3] ;
   wire \mult_21_3/FS_1/PG_int[0][3][0] ;
   wire \mult_21_3/FS_1/PG_int[0][3][1] ;
   wire \mult_21_3/A2[7] ;
   wire \mult_21_3/A2[8] ;
   wire \mult_21_3/A2[9] ;
   wire \mult_21_3/A2[10] ;
   wire \mult_21_3/A2[11] ;
   wire \mult_21_3/A2[12] ;
   wire \mult_21_3/A2[13] ;
   wire \mult_21_3/A1[0] ;
   wire \mult_21_3/A1[1] ;
   wire \mult_21_3/A1[2] ;
   wire \mult_21_3/A1[3] ;
   wire \mult_21_3/A1[4] ;
   wire \mult_21_3/A1[5] ;
   wire \mult_21_3/A1[6] ;
   wire \mult_21_3/A1[7] ;
   wire \mult_21_3/A1[8] ;
   wire \mult_21_3/A1[9] ;
   wire \mult_21_3/A1[10] ;
   wire \mult_21_3/A1[11] ;
   wire \mult_21_3/A1[12] ;
   wire \mult_21_3/ab[0][1] ;
   wire \mult_21_3/ab[0][2] ;
   wire \mult_21_3/ab[0][3] ;
   wire \mult_21_3/ab[0][4] ;
   wire \mult_21_3/ab[0][5] ;
   wire \mult_21_3/ab[0][6] ;
   wire \mult_21_3/ab[0][7] ;
   wire \mult_21_3/ab[1][0] ;
   wire \mult_21_3/ab[1][1] ;
   wire \mult_21_3/ab[1][2] ;
   wire \mult_21_3/ab[1][3] ;
   wire \mult_21_3/ab[1][4] ;
   wire \mult_21_3/ab[1][5] ;
   wire \mult_21_3/ab[1][6] ;
   wire \mult_21_3/ab[1][7] ;
   wire \mult_21_3/ab[2][0] ;
   wire \mult_21_3/ab[2][1] ;
   wire \mult_21_3/ab[2][2] ;
   wire \mult_21_3/ab[2][3] ;
   wire \mult_21_3/ab[2][4] ;
   wire \mult_21_3/ab[2][5] ;
   wire \mult_21_3/ab[2][6] ;
   wire \mult_21_3/ab[2][7] ;
   wire \mult_21_3/ab[3][0] ;
   wire \mult_21_3/ab[3][1] ;
   wire \mult_21_3/ab[3][2] ;
   wire \mult_21_3/ab[3][3] ;
   wire \mult_21_3/ab[3][4] ;
   wire \mult_21_3/ab[3][5] ;
   wire \mult_21_3/ab[3][6] ;
   wire \mult_21_3/ab[3][7] ;
   wire \mult_21_3/ab[4][0] ;
   wire \mult_21_3/ab[4][1] ;
   wire \mult_21_3/ab[4][2] ;
   wire \mult_21_3/ab[4][3] ;
   wire \mult_21_3/ab[4][4] ;
   wire \mult_21_3/ab[4][5] ;
   wire \mult_21_3/ab[4][6] ;
   wire \mult_21_3/ab[4][7] ;
   wire \mult_21_3/ab[5][0] ;
   wire \mult_21_3/ab[5][1] ;
   wire \mult_21_3/ab[5][2] ;
   wire \mult_21_3/ab[5][3] ;
   wire \mult_21_3/ab[5][4] ;
   wire \mult_21_3/ab[5][5] ;
   wire \mult_21_3/ab[5][6] ;
   wire \mult_21_3/ab[5][7] ;
   wire \mult_21_3/ab[6][0] ;
   wire \mult_21_3/ab[6][1] ;
   wire \mult_21_3/ab[6][2] ;
   wire \mult_21_3/ab[6][3] ;
   wire \mult_21_3/ab[6][4] ;
   wire \mult_21_3/ab[6][5] ;
   wire \mult_21_3/ab[6][6] ;
   wire \mult_21_3/ab[6][7] ;
   wire \mult_21_3/ab[7][0] ;
   wire \mult_21_3/ab[7][1] ;
   wire \mult_21_3/ab[7][2] ;
   wire \mult_21_3/ab[7][3] ;
   wire \mult_21_3/ab[7][4] ;
   wire \mult_21_3/ab[7][5] ;
   wire \mult_21_3/ab[7][6] ;
   wire \mult_21_3/ab[7][7] ;
   wire \mult_21_3/B_not[7] ;
   wire \mult_21_3/A_not[7] ;
   wire \mult_21_2/FS_1/C[1][2][0] ;
   wire \mult_21_2/FS_1/C[1][2][1] ;
   wire \mult_21_2/FS_1/C[1][2][2] ;
   wire \mult_21_2/FS_1/C[1][2][3] ;
   wire \mult_21_2/FS_1/C[1][3][0] ;
   wire \mult_21_2/FS_1/C[1][3][1] ;
   wire \mult_21_2/FS_1/P[0][0][1] ;
   wire \mult_21_2/FS_1/P[0][0][2] ;
   wire \mult_21_2/FS_1/P[0][0][3] ;
   wire \mult_21_2/FS_1/P[0][1][1] ;
   wire \mult_21_2/FS_1/P[0][1][2] ;
   wire \mult_21_2/FS_1/P[0][1][3] ;
   wire \mult_21_2/FS_1/P[0][2][1] ;
   wire \mult_21_2/FS_1/P[0][2][2] ;
   wire \mult_21_2/FS_1/P[0][2][3] ;
   wire \mult_21_2/FS_1/P[0][3][1] ;
   wire \mult_21_2/FS_1/TEMP_P[0][0][0] ;
   wire \mult_21_2/FS_1/TEMP_P[0][1][0] ;
   wire \mult_21_2/FS_1/TEMP_P[0][2][0] ;
   wire \mult_21_2/FS_1/TEMP_P[0][2][1] ;
   wire \mult_21_2/FS_1/TEMP_P[0][2][2] ;
   wire \mult_21_2/FS_1/TEMP_P[0][3][0] ;
   wire \mult_21_2/FS_1/G[1][0][1] ;
   wire \mult_21_2/FS_1/G[1][0][2] ;
   wire \mult_21_2/FS_1/TEMP_G[0][2][1] ;
   wire \mult_21_2/FS_1/TEMP_G[0][2][2] ;
   wire \mult_21_2/FS_1/G_n_int[0][1][3] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][0] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][1] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][2] ;
   wire \mult_21_2/FS_1/G_n_int[0][2][3] ;
   wire \mult_21_2/FS_1/G_n_int[0][3][0] ;
   wire \mult_21_2/FS_1/PG_int[0][2][0] ;
   wire \mult_21_2/FS_1/PG_int[0][2][1] ;
   wire \mult_21_2/FS_1/PG_int[0][2][2] ;
   wire \mult_21_2/FS_1/PG_int[0][2][3] ;
   wire \mult_21_2/FS_1/PG_int[0][3][0] ;
   wire \mult_21_2/FS_1/PG_int[0][3][1] ;
   wire \mult_21_2/A2[7] ;
   wire \mult_21_2/A2[8] ;
   wire \mult_21_2/A2[9] ;
   wire \mult_21_2/A2[10] ;
   wire \mult_21_2/A2[11] ;
   wire \mult_21_2/A2[12] ;
   wire \mult_21_2/A2[13] ;
   wire \mult_21_2/A1[0] ;
   wire \mult_21_2/A1[1] ;
   wire \mult_21_2/A1[2] ;
   wire \mult_21_2/A1[3] ;
   wire \mult_21_2/A1[4] ;
   wire \mult_21_2/A1[5] ;
   wire \mult_21_2/A1[6] ;
   wire \mult_21_2/A1[7] ;
   wire \mult_21_2/A1[8] ;
   wire \mult_21_2/A1[9] ;
   wire \mult_21_2/A1[10] ;
   wire \mult_21_2/A1[11] ;
   wire \mult_21_2/A1[12] ;
   wire \mult_21_2/ab[0][1] ;
   wire \mult_21_2/ab[0][2] ;
   wire \mult_21_2/ab[0][3] ;
   wire \mult_21_2/ab[0][4] ;
   wire \mult_21_2/ab[0][5] ;
   wire \mult_21_2/ab[0][6] ;
   wire \mult_21_2/ab[0][7] ;
   wire \mult_21_2/ab[1][0] ;
   wire \mult_21_2/ab[1][1] ;
   wire \mult_21_2/ab[1][2] ;
   wire \mult_21_2/ab[1][3] ;
   wire \mult_21_2/ab[1][4] ;
   wire \mult_21_2/ab[1][5] ;
   wire \mult_21_2/ab[1][6] ;
   wire \mult_21_2/ab[1][7] ;
   wire \mult_21_2/ab[2][0] ;
   wire \mult_21_2/ab[2][1] ;
   wire \mult_21_2/ab[2][2] ;
   wire \mult_21_2/ab[2][3] ;
   wire \mult_21_2/ab[2][4] ;
   wire \mult_21_2/ab[2][5] ;
   wire \mult_21_2/ab[2][6] ;
   wire \mult_21_2/ab[2][7] ;
   wire \mult_21_2/ab[3][0] ;
   wire \mult_21_2/ab[3][1] ;
   wire \mult_21_2/ab[3][2] ;
   wire \mult_21_2/ab[3][3] ;
   wire \mult_21_2/ab[3][4] ;
   wire \mult_21_2/ab[3][5] ;
   wire \mult_21_2/ab[3][6] ;
   wire \mult_21_2/ab[3][7] ;
   wire \mult_21_2/ab[4][0] ;
   wire \mult_21_2/ab[4][1] ;
   wire \mult_21_2/ab[4][2] ;
   wire \mult_21_2/ab[4][3] ;
   wire \mult_21_2/ab[4][4] ;
   wire \mult_21_2/ab[4][5] ;
   wire \mult_21_2/ab[4][6] ;
   wire \mult_21_2/ab[4][7] ;
   wire \mult_21_2/ab[5][0] ;
   wire \mult_21_2/ab[5][1] ;
   wire \mult_21_2/ab[5][2] ;
   wire \mult_21_2/ab[5][3] ;
   wire \mult_21_2/ab[5][4] ;
   wire \mult_21_2/ab[5][5] ;
   wire \mult_21_2/ab[5][6] ;
   wire \mult_21_2/ab[5][7] ;
   wire \mult_21_2/ab[6][0] ;
   wire \mult_21_2/ab[6][1] ;
   wire \mult_21_2/ab[6][2] ;
   wire \mult_21_2/ab[6][3] ;
   wire \mult_21_2/ab[6][4] ;
   wire \mult_21_2/ab[6][5] ;
   wire \mult_21_2/ab[6][6] ;
   wire \mult_21_2/ab[6][7] ;
   wire \mult_21_2/ab[7][0] ;
   wire \mult_21_2/ab[7][1] ;
   wire \mult_21_2/ab[7][2] ;
   wire \mult_21_2/ab[7][3] ;
   wire \mult_21_2/ab[7][4] ;
   wire \mult_21_2/ab[7][5] ;
   wire \mult_21_2/ab[7][6] ;
   wire \mult_21_2/ab[7][7] ;
   wire \mult_21_2/B_not[7] ;
   wire \mult_21_2/A_not[7] ;
   wire \mult_21/FS_1/C[1][2][0] ;
   wire \mult_21/FS_1/C[1][2][1] ;
   wire \mult_21/FS_1/C[1][2][2] ;
   wire \mult_21/FS_1/C[1][2][3] ;
   wire \mult_21/FS_1/C[1][3][0] ;
   wire \mult_21/FS_1/C[1][3][1] ;
   wire \mult_21/FS_1/P[0][0][1] ;
   wire \mult_21/FS_1/P[0][0][2] ;
   wire \mult_21/FS_1/P[0][0][3] ;
   wire \mult_21/FS_1/P[0][1][1] ;
   wire \mult_21/FS_1/P[0][1][2] ;
   wire \mult_21/FS_1/P[0][1][3] ;
   wire \mult_21/FS_1/P[0][2][1] ;
   wire \mult_21/FS_1/P[0][2][2] ;
   wire \mult_21/FS_1/P[0][2][3] ;
   wire \mult_21/FS_1/P[0][3][1] ;
   wire \mult_21/FS_1/TEMP_P[0][0][0] ;
   wire \mult_21/FS_1/TEMP_P[0][1][0] ;
   wire \mult_21/FS_1/TEMP_P[0][2][0] ;
   wire \mult_21/FS_1/TEMP_P[0][2][1] ;
   wire \mult_21/FS_1/TEMP_P[0][2][2] ;
   wire \mult_21/FS_1/TEMP_P[0][3][0] ;
   wire \mult_21/FS_1/G[1][0][1] ;
   wire \mult_21/FS_1/G[1][0][2] ;
   wire \mult_21/FS_1/TEMP_G[0][2][1] ;
   wire \mult_21/FS_1/TEMP_G[0][2][2] ;
   wire \mult_21/FS_1/G_n_int[0][1][3] ;
   wire \mult_21/FS_1/G_n_int[0][2][0] ;
   wire \mult_21/FS_1/G_n_int[0][2][1] ;
   wire \mult_21/FS_1/G_n_int[0][2][2] ;
   wire \mult_21/FS_1/G_n_int[0][2][3] ;
   wire \mult_21/FS_1/G_n_int[0][3][0] ;
   wire \mult_21/FS_1/PG_int[0][2][0] ;
   wire \mult_21/FS_1/PG_int[0][2][1] ;
   wire \mult_21/FS_1/PG_int[0][2][2] ;
   wire \mult_21/FS_1/PG_int[0][2][3] ;
   wire \mult_21/FS_1/PG_int[0][3][0] ;
   wire \mult_21/FS_1/PG_int[0][3][1] ;
   wire \mult_21/A2[7] ;
   wire \mult_21/A2[8] ;
   wire \mult_21/A2[9] ;
   wire \mult_21/A2[10] ;
   wire \mult_21/A2[11] ;
   wire \mult_21/A2[12] ;
   wire \mult_21/A2[13] ;
   wire \mult_21/A1[0] ;
   wire \mult_21/A1[1] ;
   wire \mult_21/A1[2] ;
   wire \mult_21/A1[3] ;
   wire \mult_21/A1[4] ;
   wire \mult_21/A1[5] ;
   wire \mult_21/A1[6] ;
   wire \mult_21/A1[7] ;
   wire \mult_21/A1[8] ;
   wire \mult_21/A1[9] ;
   wire \mult_21/A1[10] ;
   wire \mult_21/A1[11] ;
   wire \mult_21/A1[12] ;
   wire \mult_21/ab[0][1] ;
   wire \mult_21/ab[0][2] ;
   wire \mult_21/ab[0][3] ;
   wire \mult_21/ab[0][4] ;
   wire \mult_21/ab[0][5] ;
   wire \mult_21/ab[0][6] ;
   wire \mult_21/ab[0][7] ;
   wire \mult_21/ab[1][0] ;
   wire \mult_21/ab[1][1] ;
   wire \mult_21/ab[1][2] ;
   wire \mult_21/ab[1][3] ;
   wire \mult_21/ab[1][4] ;
   wire \mult_21/ab[1][5] ;
   wire \mult_21/ab[1][6] ;
   wire \mult_21/ab[1][7] ;
   wire \mult_21/ab[2][0] ;
   wire \mult_21/ab[2][1] ;
   wire \mult_21/ab[2][2] ;
   wire \mult_21/ab[2][3] ;
   wire \mult_21/ab[2][4] ;
   wire \mult_21/ab[2][5] ;
   wire \mult_21/ab[2][6] ;
   wire \mult_21/ab[2][7] ;
   wire \mult_21/ab[3][0] ;
   wire \mult_21/ab[3][1] ;
   wire \mult_21/ab[3][2] ;
   wire \mult_21/ab[3][3] ;
   wire \mult_21/ab[3][4] ;
   wire \mult_21/ab[3][5] ;
   wire \mult_21/ab[3][6] ;
   wire \mult_21/ab[3][7] ;
   wire \mult_21/ab[4][0] ;
   wire \mult_21/ab[4][1] ;
   wire \mult_21/ab[4][2] ;
   wire \mult_21/ab[4][3] ;
   wire \mult_21/ab[4][4] ;
   wire \mult_21/ab[4][5] ;
   wire \mult_21/ab[4][6] ;
   wire \mult_21/ab[4][7] ;
   wire \mult_21/ab[5][0] ;
   wire \mult_21/ab[5][1] ;
   wire \mult_21/ab[5][2] ;
   wire \mult_21/ab[5][3] ;
   wire \mult_21/ab[5][4] ;
   wire \mult_21/ab[5][5] ;
   wire \mult_21/ab[5][6] ;
   wire \mult_21/ab[5][7] ;
   wire \mult_21/ab[6][0] ;
   wire \mult_21/ab[6][1] ;
   wire \mult_21/ab[6][2] ;
   wire \mult_21/ab[6][3] ;
   wire \mult_21/ab[6][4] ;
   wire \mult_21/ab[6][5] ;
   wire \mult_21/ab[6][6] ;
   wire \mult_21/ab[6][7] ;
   wire \mult_21/ab[7][0] ;
   wire \mult_21/ab[7][1] ;
   wire \mult_21/ab[7][2] ;
   wire \mult_21/ab[7][3] ;
   wire \mult_21/ab[7][4] ;
   wire \mult_21/ab[7][5] ;
   wire \mult_21/ab[7][6] ;
   wire \mult_21/ab[7][7] ;
   wire \mult_21/B_not[7] ;
   wire \mult_21/A_not[7] ;
   wire \mult_20_3/FS_1/C[1][2][0] ;
   wire \mult_20_3/FS_1/C[1][2][1] ;
   wire \mult_20_3/FS_1/C[1][2][2] ;
   wire \mult_20_3/FS_1/C[1][2][3] ;
   wire \mult_20_3/FS_1/C[1][3][0] ;
   wire \mult_20_3/FS_1/C[1][3][1] ;
   wire \mult_20_3/FS_1/P[0][0][1] ;
   wire \mult_20_3/FS_1/P[0][0][2] ;
   wire \mult_20_3/FS_1/P[0][0][3] ;
   wire \mult_20_3/FS_1/P[0][1][1] ;
   wire \mult_20_3/FS_1/P[0][1][2] ;
   wire \mult_20_3/FS_1/P[0][1][3] ;
   wire \mult_20_3/FS_1/P[0][2][1] ;
   wire \mult_20_3/FS_1/P[0][2][2] ;
   wire \mult_20_3/FS_1/P[0][2][3] ;
   wire \mult_20_3/FS_1/P[0][3][1] ;
   wire \mult_20_3/FS_1/TEMP_P[0][0][0] ;
   wire \mult_20_3/FS_1/TEMP_P[0][1][0] ;
   wire \mult_20_3/FS_1/TEMP_P[0][2][0] ;
   wire \mult_20_3/FS_1/TEMP_P[0][2][1] ;
   wire \mult_20_3/FS_1/TEMP_P[0][2][2] ;
   wire \mult_20_3/FS_1/TEMP_P[0][3][0] ;
   wire \mult_20_3/FS_1/G[1][0][1] ;
   wire \mult_20_3/FS_1/G[1][0][2] ;
   wire \mult_20_3/FS_1/TEMP_G[0][2][1] ;
   wire \mult_20_3/FS_1/TEMP_G[0][2][2] ;
   wire \mult_20_3/FS_1/G_n_int[0][1][3] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][0] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][1] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][2] ;
   wire \mult_20_3/FS_1/G_n_int[0][2][3] ;
   wire \mult_20_3/FS_1/G_n_int[0][3][0] ;
   wire \mult_20_3/FS_1/PG_int[0][2][0] ;
   wire \mult_20_3/FS_1/PG_int[0][2][1] ;
   wire \mult_20_3/FS_1/PG_int[0][2][2] ;
   wire \mult_20_3/FS_1/PG_int[0][2][3] ;
   wire \mult_20_3/FS_1/PG_int[0][3][0] ;
   wire \mult_20_3/FS_1/PG_int[0][3][1] ;
   wire \mult_20_3/A2[7] ;
   wire \mult_20_3/A2[8] ;
   wire \mult_20_3/A2[9] ;
   wire \mult_20_3/A2[10] ;
   wire \mult_20_3/A2[11] ;
   wire \mult_20_3/A2[12] ;
   wire \mult_20_3/A2[13] ;
   wire \mult_20_3/A1[0] ;
   wire \mult_20_3/A1[1] ;
   wire \mult_20_3/A1[2] ;
   wire \mult_20_3/A1[3] ;
   wire \mult_20_3/A1[4] ;
   wire \mult_20_3/A1[5] ;
   wire \mult_20_3/A1[6] ;
   wire \mult_20_3/A1[7] ;
   wire \mult_20_3/A1[8] ;
   wire \mult_20_3/A1[9] ;
   wire \mult_20_3/A1[10] ;
   wire \mult_20_3/A1[11] ;
   wire \mult_20_3/A1[12] ;
   wire \mult_20_3/ab[0][1] ;
   wire \mult_20_3/ab[0][2] ;
   wire \mult_20_3/ab[0][3] ;
   wire \mult_20_3/ab[0][4] ;
   wire \mult_20_3/ab[0][5] ;
   wire \mult_20_3/ab[0][6] ;
   wire \mult_20_3/ab[0][7] ;
   wire \mult_20_3/ab[1][0] ;
   wire \mult_20_3/ab[1][1] ;
   wire \mult_20_3/ab[1][2] ;
   wire \mult_20_3/ab[1][3] ;
   wire \mult_20_3/ab[1][4] ;
   wire \mult_20_3/ab[1][5] ;
   wire \mult_20_3/ab[1][6] ;
   wire \mult_20_3/ab[1][7] ;
   wire \mult_20_3/ab[2][0] ;
   wire \mult_20_3/ab[2][1] ;
   wire \mult_20_3/ab[2][2] ;
   wire \mult_20_3/ab[2][3] ;
   wire \mult_20_3/ab[2][4] ;
   wire \mult_20_3/ab[2][5] ;
   wire \mult_20_3/ab[2][6] ;
   wire \mult_20_3/ab[2][7] ;
   wire \mult_20_3/ab[3][0] ;
   wire \mult_20_3/ab[3][1] ;
   wire \mult_20_3/ab[3][2] ;
   wire \mult_20_3/ab[3][3] ;
   wire \mult_20_3/ab[3][4] ;
   wire \mult_20_3/ab[3][5] ;
   wire \mult_20_3/ab[3][6] ;
   wire \mult_20_3/ab[3][7] ;
   wire \mult_20_3/ab[4][0] ;
   wire \mult_20_3/ab[4][1] ;
   wire \mult_20_3/ab[4][2] ;
   wire \mult_20_3/ab[4][3] ;
   wire \mult_20_3/ab[4][4] ;
   wire \mult_20_3/ab[4][5] ;
   wire \mult_20_3/ab[4][6] ;
   wire \mult_20_3/ab[4][7] ;
   wire \mult_20_3/ab[5][0] ;
   wire \mult_20_3/ab[5][1] ;
   wire \mult_20_3/ab[5][2] ;
   wire \mult_20_3/ab[5][3] ;
   wire \mult_20_3/ab[5][4] ;
   wire \mult_20_3/ab[5][5] ;
   wire \mult_20_3/ab[5][6] ;
   wire \mult_20_3/ab[5][7] ;
   wire \mult_20_3/ab[6][0] ;
   wire \mult_20_3/ab[6][1] ;
   wire \mult_20_3/ab[6][2] ;
   wire \mult_20_3/ab[6][3] ;
   wire \mult_20_3/ab[6][4] ;
   wire \mult_20_3/ab[6][5] ;
   wire \mult_20_3/ab[6][6] ;
   wire \mult_20_3/ab[6][7] ;
   wire \mult_20_3/ab[7][0] ;
   wire \mult_20_3/ab[7][1] ;
   wire \mult_20_3/ab[7][2] ;
   wire \mult_20_3/ab[7][3] ;
   wire \mult_20_3/ab[7][4] ;
   wire \mult_20_3/ab[7][5] ;
   wire \mult_20_3/ab[7][6] ;
   wire \mult_20_3/ab[7][7] ;
   wire \mult_20_3/B_not[7] ;
   wire \mult_20_3/A_not[7] ;
   wire \mult_20_2/FS_1/C[1][2][0] ;
   wire \mult_20_2/FS_1/C[1][2][1] ;
   wire \mult_20_2/FS_1/C[1][2][2] ;
   wire \mult_20_2/FS_1/C[1][2][3] ;
   wire \mult_20_2/FS_1/C[1][3][0] ;
   wire \mult_20_2/FS_1/C[1][3][1] ;
   wire \mult_20_2/FS_1/P[0][0][1] ;
   wire \mult_20_2/FS_1/P[0][0][2] ;
   wire \mult_20_2/FS_1/P[0][0][3] ;
   wire \mult_20_2/FS_1/P[0][1][1] ;
   wire \mult_20_2/FS_1/P[0][1][2] ;
   wire \mult_20_2/FS_1/P[0][1][3] ;
   wire \mult_20_2/FS_1/P[0][2][1] ;
   wire \mult_20_2/FS_1/P[0][2][2] ;
   wire \mult_20_2/FS_1/P[0][2][3] ;
   wire \mult_20_2/FS_1/P[0][3][1] ;
   wire \mult_20_2/FS_1/TEMP_P[0][0][0] ;
   wire \mult_20_2/FS_1/TEMP_P[0][1][0] ;
   wire \mult_20_2/FS_1/TEMP_P[0][2][0] ;
   wire \mult_20_2/FS_1/TEMP_P[0][2][1] ;
   wire \mult_20_2/FS_1/TEMP_P[0][2][2] ;
   wire \mult_20_2/FS_1/TEMP_P[0][3][0] ;
   wire \mult_20_2/FS_1/G[1][0][1] ;
   wire \mult_20_2/FS_1/G[1][0][2] ;
   wire \mult_20_2/FS_1/TEMP_G[0][2][1] ;
   wire \mult_20_2/FS_1/TEMP_G[0][2][2] ;
   wire \mult_20_2/FS_1/G_n_int[0][1][3] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][0] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][1] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][2] ;
   wire \mult_20_2/FS_1/G_n_int[0][2][3] ;
   wire \mult_20_2/FS_1/G_n_int[0][3][0] ;
   wire \mult_20_2/FS_1/PG_int[0][2][0] ;
   wire \mult_20_2/FS_1/PG_int[0][2][1] ;
   wire \mult_20_2/FS_1/PG_int[0][2][2] ;
   wire \mult_20_2/FS_1/PG_int[0][2][3] ;
   wire \mult_20_2/FS_1/PG_int[0][3][0] ;
   wire \mult_20_2/FS_1/PG_int[0][3][1] ;
   wire \mult_20_2/A2[7] ;
   wire \mult_20_2/A2[8] ;
   wire \mult_20_2/A2[9] ;
   wire \mult_20_2/A2[10] ;
   wire \mult_20_2/A2[11] ;
   wire \mult_20_2/A2[12] ;
   wire \mult_20_2/A2[13] ;
   wire \mult_20_2/A1[0] ;
   wire \mult_20_2/A1[1] ;
   wire \mult_20_2/A1[2] ;
   wire \mult_20_2/A1[3] ;
   wire \mult_20_2/A1[4] ;
   wire \mult_20_2/A1[5] ;
   wire \mult_20_2/A1[6] ;
   wire \mult_20_2/A1[7] ;
   wire \mult_20_2/A1[8] ;
   wire \mult_20_2/A1[9] ;
   wire \mult_20_2/A1[10] ;
   wire \mult_20_2/A1[11] ;
   wire \mult_20_2/A1[12] ;
   wire \mult_20_2/ab[0][1] ;
   wire \mult_20_2/ab[0][2] ;
   wire \mult_20_2/ab[0][3] ;
   wire \mult_20_2/ab[0][4] ;
   wire \mult_20_2/ab[0][5] ;
   wire \mult_20_2/ab[0][6] ;
   wire \mult_20_2/ab[0][7] ;
   wire \mult_20_2/ab[1][0] ;
   wire \mult_20_2/ab[1][1] ;
   wire \mult_20_2/ab[1][2] ;
   wire \mult_20_2/ab[1][3] ;
   wire \mult_20_2/ab[1][4] ;
   wire \mult_20_2/ab[1][5] ;
   wire \mult_20_2/ab[1][6] ;
   wire \mult_20_2/ab[1][7] ;
   wire \mult_20_2/ab[2][0] ;
   wire \mult_20_2/ab[2][1] ;
   wire \mult_20_2/ab[2][2] ;
   wire \mult_20_2/ab[2][3] ;
   wire \mult_20_2/ab[2][4] ;
   wire \mult_20_2/ab[2][5] ;
   wire \mult_20_2/ab[2][6] ;
   wire \mult_20_2/ab[2][7] ;
   wire \mult_20_2/ab[3][0] ;
   wire \mult_20_2/ab[3][1] ;
   wire \mult_20_2/ab[3][2] ;
   wire \mult_20_2/ab[3][3] ;
   wire \mult_20_2/ab[3][4] ;
   wire \mult_20_2/ab[3][5] ;
   wire \mult_20_2/ab[3][6] ;
   wire \mult_20_2/ab[3][7] ;
   wire \mult_20_2/ab[4][0] ;
   wire \mult_20_2/ab[4][1] ;
   wire \mult_20_2/ab[4][2] ;
   wire \mult_20_2/ab[4][3] ;
   wire \mult_20_2/ab[4][4] ;
   wire \mult_20_2/ab[4][5] ;
   wire \mult_20_2/ab[4][6] ;
   wire \mult_20_2/ab[4][7] ;
   wire \mult_20_2/ab[5][0] ;
   wire \mult_20_2/ab[5][1] ;
   wire \mult_20_2/ab[5][2] ;
   wire \mult_20_2/ab[5][3] ;
   wire \mult_20_2/ab[5][4] ;
   wire \mult_20_2/ab[5][5] ;
   wire \mult_20_2/ab[5][6] ;
   wire \mult_20_2/ab[5][7] ;
   wire \mult_20_2/ab[6][0] ;
   wire \mult_20_2/ab[6][1] ;
   wire \mult_20_2/ab[6][2] ;
   wire \mult_20_2/ab[6][3] ;
   wire \mult_20_2/ab[6][4] ;
   wire \mult_20_2/ab[6][5] ;
   wire \mult_20_2/ab[6][6] ;
   wire \mult_20_2/ab[6][7] ;
   wire \mult_20_2/ab[7][0] ;
   wire \mult_20_2/ab[7][1] ;
   wire \mult_20_2/ab[7][2] ;
   wire \mult_20_2/ab[7][3] ;
   wire \mult_20_2/ab[7][4] ;
   wire \mult_20_2/ab[7][5] ;
   wire \mult_20_2/ab[7][6] ;
   wire \mult_20_2/ab[7][7] ;
   wire \mult_20_2/B_not[7] ;
   wire \mult_20_2/A_not[7] ;
   wire \mult_20/FS_1/C[1][2][0] ;
   wire \mult_20/FS_1/C[1][2][1] ;
   wire \mult_20/FS_1/C[1][2][2] ;
   wire \mult_20/FS_1/C[1][2][3] ;
   wire \mult_20/FS_1/C[1][3][0] ;
   wire \mult_20/FS_1/C[1][3][1] ;
   wire \mult_20/FS_1/P[0][0][1] ;
   wire \mult_20/FS_1/P[0][0][2] ;
   wire \mult_20/FS_1/P[0][0][3] ;
   wire \mult_20/FS_1/P[0][1][1] ;
   wire \mult_20/FS_1/P[0][1][2] ;
   wire \mult_20/FS_1/P[0][1][3] ;
   wire \mult_20/FS_1/P[0][2][1] ;
   wire \mult_20/FS_1/P[0][2][2] ;
   wire \mult_20/FS_1/P[0][2][3] ;
   wire \mult_20/FS_1/P[0][3][1] ;
   wire \mult_20/FS_1/TEMP_P[0][0][0] ;
   wire \mult_20/FS_1/TEMP_P[0][1][0] ;
   wire \mult_20/FS_1/TEMP_P[0][2][0] ;
   wire \mult_20/FS_1/TEMP_P[0][2][1] ;
   wire \mult_20/FS_1/TEMP_P[0][2][2] ;
   wire \mult_20/FS_1/TEMP_P[0][3][0] ;
   wire \mult_20/FS_1/G[1][0][1] ;
   wire \mult_20/FS_1/G[1][0][2] ;
   wire \mult_20/FS_1/TEMP_G[0][2][1] ;
   wire \mult_20/FS_1/TEMP_G[0][2][2] ;
   wire \mult_20/FS_1/G_n_int[0][1][3] ;
   wire \mult_20/FS_1/G_n_int[0][2][0] ;
   wire \mult_20/FS_1/G_n_int[0][2][1] ;
   wire \mult_20/FS_1/G_n_int[0][2][2] ;
   wire \mult_20/FS_1/G_n_int[0][2][3] ;
   wire \mult_20/FS_1/G_n_int[0][3][0] ;
   wire \mult_20/FS_1/PG_int[0][2][0] ;
   wire \mult_20/FS_1/PG_int[0][2][1] ;
   wire \mult_20/FS_1/PG_int[0][2][2] ;
   wire \mult_20/FS_1/PG_int[0][2][3] ;
   wire \mult_20/FS_1/PG_int[0][3][0] ;
   wire \mult_20/FS_1/PG_int[0][3][1] ;
   wire \mult_20/A2[7] ;
   wire \mult_20/A2[8] ;
   wire \mult_20/A2[9] ;
   wire \mult_20/A2[10] ;
   wire \mult_20/A2[11] ;
   wire \mult_20/A2[12] ;
   wire \mult_20/A2[13] ;
   wire \mult_20/A1[0] ;
   wire \mult_20/A1[1] ;
   wire \mult_20/A1[2] ;
   wire \mult_20/A1[3] ;
   wire \mult_20/A1[4] ;
   wire \mult_20/A1[5] ;
   wire \mult_20/A1[6] ;
   wire \mult_20/A1[7] ;
   wire \mult_20/A1[8] ;
   wire \mult_20/A1[9] ;
   wire \mult_20/A1[10] ;
   wire \mult_20/A1[11] ;
   wire \mult_20/A1[12] ;
   wire \mult_20/ab[0][1] ;
   wire \mult_20/ab[0][2] ;
   wire \mult_20/ab[0][3] ;
   wire \mult_20/ab[0][4] ;
   wire \mult_20/ab[0][5] ;
   wire \mult_20/ab[0][6] ;
   wire \mult_20/ab[0][7] ;
   wire \mult_20/ab[1][0] ;
   wire \mult_20/ab[1][1] ;
   wire \mult_20/ab[1][2] ;
   wire \mult_20/ab[1][3] ;
   wire \mult_20/ab[1][4] ;
   wire \mult_20/ab[1][5] ;
   wire \mult_20/ab[1][6] ;
   wire \mult_20/ab[1][7] ;
   wire \mult_20/ab[2][0] ;
   wire \mult_20/ab[2][1] ;
   wire \mult_20/ab[2][2] ;
   wire \mult_20/ab[2][3] ;
   wire \mult_20/ab[2][4] ;
   wire \mult_20/ab[2][5] ;
   wire \mult_20/ab[2][6] ;
   wire \mult_20/ab[2][7] ;
   wire \mult_20/ab[3][0] ;
   wire \mult_20/ab[3][1] ;
   wire \mult_20/ab[3][2] ;
   wire \mult_20/ab[3][3] ;
   wire \mult_20/ab[3][4] ;
   wire \mult_20/ab[3][5] ;
   wire \mult_20/ab[3][6] ;
   wire \mult_20/ab[3][7] ;
   wire \mult_20/ab[4][0] ;
   wire \mult_20/ab[4][1] ;
   wire \mult_20/ab[4][2] ;
   wire \mult_20/ab[4][3] ;
   wire \mult_20/ab[4][4] ;
   wire \mult_20/ab[4][5] ;
   wire \mult_20/ab[4][6] ;
   wire \mult_20/ab[4][7] ;
   wire \mult_20/ab[5][0] ;
   wire \mult_20/ab[5][1] ;
   wire \mult_20/ab[5][2] ;
   wire \mult_20/ab[5][3] ;
   wire \mult_20/ab[5][4] ;
   wire \mult_20/ab[5][5] ;
   wire \mult_20/ab[5][6] ;
   wire \mult_20/ab[5][7] ;
   wire \mult_20/ab[6][0] ;
   wire \mult_20/ab[6][1] ;
   wire \mult_20/ab[6][2] ;
   wire \mult_20/ab[6][3] ;
   wire \mult_20/ab[6][4] ;
   wire \mult_20/ab[6][5] ;
   wire \mult_20/ab[6][6] ;
   wire \mult_20/ab[6][7] ;
   wire \mult_20/ab[7][0] ;
   wire \mult_20/ab[7][1] ;
   wire \mult_20/ab[7][2] ;
   wire \mult_20/ab[7][3] ;
   wire \mult_20/ab[7][4] ;
   wire \mult_20/ab[7][5] ;
   wire \mult_20/ab[7][6] ;
   wire \mult_20/ab[7][7] ;
   wire \mult_20/B_not[7] ;
   wire \mult_20/A_not[7] ;
   wire \mult_19_3/FS_1/C[1][2][0] ;
   wire \mult_19_3/FS_1/C[1][2][1] ;
   wire \mult_19_3/FS_1/C[1][2][2] ;
   wire \mult_19_3/FS_1/C[1][2][3] ;
   wire \mult_19_3/FS_1/C[1][3][0] ;
   wire \mult_19_3/FS_1/C[1][3][1] ;
   wire \mult_19_3/FS_1/P[0][0][1] ;
   wire \mult_19_3/FS_1/P[0][0][2] ;
   wire \mult_19_3/FS_1/P[0][0][3] ;
   wire \mult_19_3/FS_1/P[0][1][1] ;
   wire \mult_19_3/FS_1/P[0][1][2] ;
   wire \mult_19_3/FS_1/P[0][1][3] ;
   wire \mult_19_3/FS_1/P[0][2][1] ;
   wire \mult_19_3/FS_1/P[0][2][2] ;
   wire \mult_19_3/FS_1/P[0][2][3] ;
   wire \mult_19_3/FS_1/P[0][3][1] ;
   wire \mult_19_3/FS_1/TEMP_P[0][0][0] ;
   wire \mult_19_3/FS_1/TEMP_P[0][1][0] ;
   wire \mult_19_3/FS_1/TEMP_P[0][2][0] ;
   wire \mult_19_3/FS_1/TEMP_P[0][2][1] ;
   wire \mult_19_3/FS_1/TEMP_P[0][2][2] ;
   wire \mult_19_3/FS_1/TEMP_P[0][3][0] ;
   wire \mult_19_3/FS_1/G[1][0][1] ;
   wire \mult_19_3/FS_1/G[1][0][2] ;
   wire \mult_19_3/FS_1/TEMP_G[0][2][1] ;
   wire \mult_19_3/FS_1/TEMP_G[0][2][2] ;
   wire \mult_19_3/FS_1/G_n_int[0][1][3] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][0] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][1] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][2] ;
   wire \mult_19_3/FS_1/G_n_int[0][2][3] ;
   wire \mult_19_3/FS_1/G_n_int[0][3][0] ;
   wire \mult_19_3/FS_1/PG_int[0][2][0] ;
   wire \mult_19_3/FS_1/PG_int[0][2][1] ;
   wire \mult_19_3/FS_1/PG_int[0][2][2] ;
   wire \mult_19_3/FS_1/PG_int[0][2][3] ;
   wire \mult_19_3/FS_1/PG_int[0][3][0] ;
   wire \mult_19_3/FS_1/PG_int[0][3][1] ;
   wire \mult_19_3/A2[7] ;
   wire \mult_19_3/A2[8] ;
   wire \mult_19_3/A2[9] ;
   wire \mult_19_3/A2[10] ;
   wire \mult_19_3/A2[11] ;
   wire \mult_19_3/A2[12] ;
   wire \mult_19_3/A2[13] ;
   wire \mult_19_3/A1[0] ;
   wire \mult_19_3/A1[1] ;
   wire \mult_19_3/A1[2] ;
   wire \mult_19_3/A1[3] ;
   wire \mult_19_3/A1[4] ;
   wire \mult_19_3/A1[5] ;
   wire \mult_19_3/A1[6] ;
   wire \mult_19_3/A1[7] ;
   wire \mult_19_3/A1[8] ;
   wire \mult_19_3/A1[9] ;
   wire \mult_19_3/A1[10] ;
   wire \mult_19_3/A1[11] ;
   wire \mult_19_3/A1[12] ;
   wire \mult_19_3/ab[0][1] ;
   wire \mult_19_3/ab[0][2] ;
   wire \mult_19_3/ab[0][3] ;
   wire \mult_19_3/ab[0][4] ;
   wire \mult_19_3/ab[0][5] ;
   wire \mult_19_3/ab[0][6] ;
   wire \mult_19_3/ab[0][7] ;
   wire \mult_19_3/ab[1][0] ;
   wire \mult_19_3/ab[1][1] ;
   wire \mult_19_3/ab[1][2] ;
   wire \mult_19_3/ab[1][3] ;
   wire \mult_19_3/ab[1][4] ;
   wire \mult_19_3/ab[1][5] ;
   wire \mult_19_3/ab[1][6] ;
   wire \mult_19_3/ab[1][7] ;
   wire \mult_19_3/ab[2][0] ;
   wire \mult_19_3/ab[2][1] ;
   wire \mult_19_3/ab[2][2] ;
   wire \mult_19_3/ab[2][3] ;
   wire \mult_19_3/ab[2][4] ;
   wire \mult_19_3/ab[2][5] ;
   wire \mult_19_3/ab[2][6] ;
   wire \mult_19_3/ab[2][7] ;
   wire \mult_19_3/ab[3][0] ;
   wire \mult_19_3/ab[3][1] ;
   wire \mult_19_3/ab[3][2] ;
   wire \mult_19_3/ab[3][3] ;
   wire \mult_19_3/ab[3][4] ;
   wire \mult_19_3/ab[3][5] ;
   wire \mult_19_3/ab[3][6] ;
   wire \mult_19_3/ab[3][7] ;
   wire \mult_19_3/ab[4][0] ;
   wire \mult_19_3/ab[4][1] ;
   wire \mult_19_3/ab[4][2] ;
   wire \mult_19_3/ab[4][3] ;
   wire \mult_19_3/ab[4][4] ;
   wire \mult_19_3/ab[4][5] ;
   wire \mult_19_3/ab[4][6] ;
   wire \mult_19_3/ab[4][7] ;
   wire \mult_19_3/ab[5][0] ;
   wire \mult_19_3/ab[5][1] ;
   wire \mult_19_3/ab[5][2] ;
   wire \mult_19_3/ab[5][3] ;
   wire \mult_19_3/ab[5][4] ;
   wire \mult_19_3/ab[5][5] ;
   wire \mult_19_3/ab[5][6] ;
   wire \mult_19_3/ab[5][7] ;
   wire \mult_19_3/ab[6][0] ;
   wire \mult_19_3/ab[6][1] ;
   wire \mult_19_3/ab[6][2] ;
   wire \mult_19_3/ab[6][3] ;
   wire \mult_19_3/ab[6][4] ;
   wire \mult_19_3/ab[6][5] ;
   wire \mult_19_3/ab[6][6] ;
   wire \mult_19_3/ab[6][7] ;
   wire \mult_19_3/ab[7][0] ;
   wire \mult_19_3/ab[7][1] ;
   wire \mult_19_3/ab[7][2] ;
   wire \mult_19_3/ab[7][3] ;
   wire \mult_19_3/ab[7][4] ;
   wire \mult_19_3/ab[7][5] ;
   wire \mult_19_3/ab[7][6] ;
   wire \mult_19_3/ab[7][7] ;
   wire \mult_19_3/B_not[7] ;
   wire \mult_19_3/A_not[7] ;
   wire \mult_19_2/FS_1/C[1][2][0] ;
   wire \mult_19_2/FS_1/C[1][2][1] ;
   wire \mult_19_2/FS_1/C[1][2][2] ;
   wire \mult_19_2/FS_1/C[1][2][3] ;
   wire \mult_19_2/FS_1/C[1][3][0] ;
   wire \mult_19_2/FS_1/C[1][3][1] ;
   wire \mult_19_2/FS_1/P[0][0][1] ;
   wire \mult_19_2/FS_1/P[0][0][2] ;
   wire \mult_19_2/FS_1/P[0][0][3] ;
   wire \mult_19_2/FS_1/P[0][1][1] ;
   wire \mult_19_2/FS_1/P[0][1][2] ;
   wire \mult_19_2/FS_1/P[0][1][3] ;
   wire \mult_19_2/FS_1/P[0][2][1] ;
   wire \mult_19_2/FS_1/P[0][2][2] ;
   wire \mult_19_2/FS_1/P[0][2][3] ;
   wire \mult_19_2/FS_1/P[0][3][1] ;
   wire \mult_19_2/FS_1/TEMP_P[0][0][0] ;
   wire \mult_19_2/FS_1/TEMP_P[0][1][0] ;
   wire \mult_19_2/FS_1/TEMP_P[0][2][0] ;
   wire \mult_19_2/FS_1/TEMP_P[0][2][1] ;
   wire \mult_19_2/FS_1/TEMP_P[0][2][2] ;
   wire \mult_19_2/FS_1/TEMP_P[0][3][0] ;
   wire \mult_19_2/FS_1/G[1][0][1] ;
   wire \mult_19_2/FS_1/G[1][0][2] ;
   wire \mult_19_2/FS_1/TEMP_G[0][2][1] ;
   wire \mult_19_2/FS_1/TEMP_G[0][2][2] ;
   wire \mult_19_2/FS_1/G_n_int[0][1][3] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][0] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][1] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][2] ;
   wire \mult_19_2/FS_1/G_n_int[0][2][3] ;
   wire \mult_19_2/FS_1/G_n_int[0][3][0] ;
   wire \mult_19_2/FS_1/PG_int[0][2][0] ;
   wire \mult_19_2/FS_1/PG_int[0][2][1] ;
   wire \mult_19_2/FS_1/PG_int[0][2][2] ;
   wire \mult_19_2/FS_1/PG_int[0][2][3] ;
   wire \mult_19_2/FS_1/PG_int[0][3][0] ;
   wire \mult_19_2/FS_1/PG_int[0][3][1] ;
   wire \mult_19_2/A2[7] ;
   wire \mult_19_2/A2[8] ;
   wire \mult_19_2/A2[9] ;
   wire \mult_19_2/A2[10] ;
   wire \mult_19_2/A2[11] ;
   wire \mult_19_2/A2[12] ;
   wire \mult_19_2/A2[13] ;
   wire \mult_19_2/A1[0] ;
   wire \mult_19_2/A1[1] ;
   wire \mult_19_2/A1[2] ;
   wire \mult_19_2/A1[3] ;
   wire \mult_19_2/A1[4] ;
   wire \mult_19_2/A1[5] ;
   wire \mult_19_2/A1[6] ;
   wire \mult_19_2/A1[7] ;
   wire \mult_19_2/A1[8] ;
   wire \mult_19_2/A1[9] ;
   wire \mult_19_2/A1[10] ;
   wire \mult_19_2/A1[11] ;
   wire \mult_19_2/A1[12] ;
   wire \mult_19_2/ab[0][1] ;
   wire \mult_19_2/ab[0][2] ;
   wire \mult_19_2/ab[0][3] ;
   wire \mult_19_2/ab[0][4] ;
   wire \mult_19_2/ab[0][5] ;
   wire \mult_19_2/ab[0][6] ;
   wire \mult_19_2/ab[0][7] ;
   wire \mult_19_2/ab[1][0] ;
   wire \mult_19_2/ab[1][1] ;
   wire \mult_19_2/ab[1][2] ;
   wire \mult_19_2/ab[1][3] ;
   wire \mult_19_2/ab[1][4] ;
   wire \mult_19_2/ab[1][5] ;
   wire \mult_19_2/ab[1][6] ;
   wire \mult_19_2/ab[1][7] ;
   wire \mult_19_2/ab[2][0] ;
   wire \mult_19_2/ab[2][1] ;
   wire \mult_19_2/ab[2][2] ;
   wire \mult_19_2/ab[2][3] ;
   wire \mult_19_2/ab[2][4] ;
   wire \mult_19_2/ab[2][5] ;
   wire \mult_19_2/ab[2][6] ;
   wire \mult_19_2/ab[2][7] ;
   wire \mult_19_2/ab[3][0] ;
   wire \mult_19_2/ab[3][1] ;
   wire \mult_19_2/ab[3][2] ;
   wire \mult_19_2/ab[3][3] ;
   wire \mult_19_2/ab[3][4] ;
   wire \mult_19_2/ab[3][5] ;
   wire \mult_19_2/ab[3][6] ;
   wire \mult_19_2/ab[3][7] ;
   wire \mult_19_2/ab[4][0] ;
   wire \mult_19_2/ab[4][1] ;
   wire \mult_19_2/ab[4][2] ;
   wire \mult_19_2/ab[4][3] ;
   wire \mult_19_2/ab[4][4] ;
   wire \mult_19_2/ab[4][5] ;
   wire \mult_19_2/ab[4][6] ;
   wire \mult_19_2/ab[4][7] ;
   wire \mult_19_2/ab[5][0] ;
   wire \mult_19_2/ab[5][1] ;
   wire \mult_19_2/ab[5][2] ;
   wire \mult_19_2/ab[5][3] ;
   wire \mult_19_2/ab[5][4] ;
   wire \mult_19_2/ab[5][5] ;
   wire \mult_19_2/ab[5][6] ;
   wire \mult_19_2/ab[5][7] ;
   wire \mult_19_2/ab[6][0] ;
   wire \mult_19_2/ab[6][1] ;
   wire \mult_19_2/ab[6][2] ;
   wire \mult_19_2/ab[6][3] ;
   wire \mult_19_2/ab[6][4] ;
   wire \mult_19_2/ab[6][5] ;
   wire \mult_19_2/ab[6][6] ;
   wire \mult_19_2/ab[6][7] ;
   wire \mult_19_2/ab[7][0] ;
   wire \mult_19_2/ab[7][1] ;
   wire \mult_19_2/ab[7][2] ;
   wire \mult_19_2/ab[7][3] ;
   wire \mult_19_2/ab[7][4] ;
   wire \mult_19_2/ab[7][5] ;
   wire \mult_19_2/ab[7][6] ;
   wire \mult_19_2/ab[7][7] ;
   wire \mult_19_2/B_not[7] ;
   wire \mult_19_2/A_not[7] ;
   wire \mult_19/FS_1/C[1][2][0] ;
   wire \mult_19/FS_1/C[1][2][1] ;
   wire \mult_19/FS_1/C[1][2][2] ;
   wire \mult_19/FS_1/C[1][2][3] ;
   wire \mult_19/FS_1/C[1][3][0] ;
   wire \mult_19/FS_1/C[1][3][1] ;
   wire \mult_19/FS_1/P[0][0][1] ;
   wire \mult_19/FS_1/P[0][0][2] ;
   wire \mult_19/FS_1/P[0][0][3] ;
   wire \mult_19/FS_1/P[0][1][1] ;
   wire \mult_19/FS_1/P[0][1][2] ;
   wire \mult_19/FS_1/P[0][1][3] ;
   wire \mult_19/FS_1/P[0][2][1] ;
   wire \mult_19/FS_1/P[0][2][2] ;
   wire \mult_19/FS_1/P[0][2][3] ;
   wire \mult_19/FS_1/P[0][3][1] ;
   wire \mult_19/FS_1/TEMP_P[0][0][0] ;
   wire \mult_19/FS_1/TEMP_P[0][1][0] ;
   wire \mult_19/FS_1/TEMP_P[0][2][0] ;
   wire \mult_19/FS_1/TEMP_P[0][2][1] ;
   wire \mult_19/FS_1/TEMP_P[0][2][2] ;
   wire \mult_19/FS_1/TEMP_P[0][3][0] ;
   wire \mult_19/FS_1/G[1][0][1] ;
   wire \mult_19/FS_1/G[1][0][2] ;
   wire \mult_19/FS_1/TEMP_G[0][2][1] ;
   wire \mult_19/FS_1/TEMP_G[0][2][2] ;
   wire \mult_19/FS_1/G_n_int[0][1][3] ;
   wire \mult_19/FS_1/G_n_int[0][2][0] ;
   wire \mult_19/FS_1/G_n_int[0][2][1] ;
   wire \mult_19/FS_1/G_n_int[0][2][2] ;
   wire \mult_19/FS_1/G_n_int[0][2][3] ;
   wire \mult_19/FS_1/G_n_int[0][3][0] ;
   wire \mult_19/FS_1/PG_int[0][2][0] ;
   wire \mult_19/FS_1/PG_int[0][2][1] ;
   wire \mult_19/FS_1/PG_int[0][2][2] ;
   wire \mult_19/FS_1/PG_int[0][2][3] ;
   wire \mult_19/FS_1/PG_int[0][3][0] ;
   wire \mult_19/FS_1/PG_int[0][3][1] ;
   wire \mult_19/A2[7] ;
   wire \mult_19/A2[8] ;
   wire \mult_19/A2[9] ;
   wire \mult_19/A2[10] ;
   wire \mult_19/A2[11] ;
   wire \mult_19/A2[12] ;
   wire \mult_19/A2[13] ;
   wire \mult_19/A1[0] ;
   wire \mult_19/A1[1] ;
   wire \mult_19/A1[2] ;
   wire \mult_19/A1[3] ;
   wire \mult_19/A1[4] ;
   wire \mult_19/A1[5] ;
   wire \mult_19/A1[6] ;
   wire \mult_19/A1[7] ;
   wire \mult_19/A1[8] ;
   wire \mult_19/A1[9] ;
   wire \mult_19/A1[10] ;
   wire \mult_19/A1[11] ;
   wire \mult_19/A1[12] ;
   wire \mult_19/ab[0][1] ;
   wire \mult_19/ab[0][2] ;
   wire \mult_19/ab[0][3] ;
   wire \mult_19/ab[0][4] ;
   wire \mult_19/ab[0][5] ;
   wire \mult_19/ab[0][6] ;
   wire \mult_19/ab[0][7] ;
   wire \mult_19/ab[1][0] ;
   wire \mult_19/ab[1][1] ;
   wire \mult_19/ab[1][2] ;
   wire \mult_19/ab[1][3] ;
   wire \mult_19/ab[1][4] ;
   wire \mult_19/ab[1][5] ;
   wire \mult_19/ab[1][6] ;
   wire \mult_19/ab[1][7] ;
   wire \mult_19/ab[2][0] ;
   wire \mult_19/ab[2][1] ;
   wire \mult_19/ab[2][2] ;
   wire \mult_19/ab[2][3] ;
   wire \mult_19/ab[2][4] ;
   wire \mult_19/ab[2][5] ;
   wire \mult_19/ab[2][6] ;
   wire \mult_19/ab[2][7] ;
   wire \mult_19/ab[3][0] ;
   wire \mult_19/ab[3][1] ;
   wire \mult_19/ab[3][2] ;
   wire \mult_19/ab[3][3] ;
   wire \mult_19/ab[3][4] ;
   wire \mult_19/ab[3][5] ;
   wire \mult_19/ab[3][6] ;
   wire \mult_19/ab[3][7] ;
   wire \mult_19/ab[4][0] ;
   wire \mult_19/ab[4][1] ;
   wire \mult_19/ab[4][2] ;
   wire \mult_19/ab[4][3] ;
   wire \mult_19/ab[4][4] ;
   wire \mult_19/ab[4][5] ;
   wire \mult_19/ab[4][6] ;
   wire \mult_19/ab[4][7] ;
   wire \mult_19/ab[5][0] ;
   wire \mult_19/ab[5][1] ;
   wire \mult_19/ab[5][2] ;
   wire \mult_19/ab[5][3] ;
   wire \mult_19/ab[5][4] ;
   wire \mult_19/ab[5][5] ;
   wire \mult_19/ab[5][6] ;
   wire \mult_19/ab[5][7] ;
   wire \mult_19/ab[6][0] ;
   wire \mult_19/ab[6][1] ;
   wire \mult_19/ab[6][2] ;
   wire \mult_19/ab[6][3] ;
   wire \mult_19/ab[6][4] ;
   wire \mult_19/ab[6][5] ;
   wire \mult_19/ab[6][6] ;
   wire \mult_19/ab[6][7] ;
   wire \mult_19/ab[7][0] ;
   wire \mult_19/ab[7][1] ;
   wire \mult_19/ab[7][2] ;
   wire \mult_19/ab[7][3] ;
   wire \mult_19/ab[7][4] ;
   wire \mult_19/ab[7][5] ;
   wire \mult_19/ab[7][6] ;
   wire \mult_19/ab[7][7] ;
   wire \mult_19/B_not[7] ;
   wire \mult_19/A_not[7] ;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3297;
   wire n3298;
   wire n3299;
   wire n3300;
   wire n3301;
   wire n3302;
   wire n3303;
   wire n3304;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire [6:0] \mult_21_3/A_notx ;
   wire [6:0] \mult_21_3/B_notx ;
   wire [6:0] \mult_21_2/A_notx ;
   wire [6:0] \mult_21_2/B_notx ;
   wire [6:0] \mult_21/A_notx ;
   wire [6:0] \mult_21/B_notx ;
   wire [6:0] \mult_20_3/A_notx ;
   wire [6:0] \mult_20_3/B_notx ;
   wire [6:0] \mult_20_2/A_notx ;
   wire [6:0] \mult_20_2/B_notx ;
   wire [6:0] \mult_20/A_notx ;
   wire [6:0] \mult_20/B_notx ;
   wire [6:0] \mult_19_3/A_notx ;
   wire [6:0] \mult_19_3/B_notx ;
   wire [6:0] \mult_19_2/A_notx ;
   wire [6:0] \mult_19_2/B_notx ;
   wire [6:0] \mult_19/A_notx ;
   wire [6:0] \mult_19/B_notx ;

   INVERTER I_0 (.IN(rst_n),
	.OUT(N0));
   DFF \result_1_reg[15]  (.D(N160),
	.CLK(n53),
	.R(N0),
	.Q(result_1[15]));
   DFF \result_1_reg[14]  (.D(N159),
	.CLK(n32),
	.R(n54),
	.Q(result_1[14]));
   DFF \result_1_reg[13]  (.D(N158),
	.CLK(n21),
	.R(n55),
	.Q(result_1[13]));
   DFF \result_1_reg[12]  (.D(N157),
	.CLK(n39),
	.R(N0),
	.Q(result_1[12]));
   DFF \result_1_reg[11]  (.D(N156),
	.CLK(n61),
	.R(n54),
	.Q(result_1[11]));
   DFF \result_1_reg[10]  (.D(N155),
	.CLK(n1),
	.R(n55),
	.Q(result_1[10]));
   DFF \result_1_reg[9]  (.D(N154),
	.CLK(n43),
	.R(N0),
	.Q(result_1[9]));
   DFF \result_1_reg[8]  (.D(N153),
	.CLK(n47),
	.R(n54),
	.Q(result_1[8]));
   DFF \result_1_reg[7]  (.D(N152),
	.CLK(n52),
	.R(n55),
	.Q(result_1[7]));
   DFF \result_1_reg[6]  (.D(N151),
	.CLK(n17),
	.R(N0),
	.Q(result_1[6]));
   DFF \result_1_reg[5]  (.D(N150),
	.CLK(n45),
	.R(n54),
	.Q(result_1[5]));
   DFF \result_1_reg[4]  (.D(N149),
	.CLK(n44),
	.R(n55),
	.Q(result_1[4]));
   DFF \result_1_reg[3]  (.D(N148),
	.CLK(n40),
	.R(N0),
	.Q(result_1[3]));
   DFF \result_1_reg[2]  (.D(N147),
	.CLK(n23),
	.R(n54),
	.Q(result_1[2]));
   DFF \result_1_reg[1]  (.D(N146),
	.CLK(n38),
	.R(n55),
	.Q(result_1[1]));
   DFF \result_1_reg[0]  (.D(N145),
	.CLK(n34),
	.R(N0),
	.Q(result_1[0]));
   DFF \result_2_reg[15]  (.D(N240),
	.CLK(n28),
	.R(n54),
	.Q(result_2[15]));
   DFF \result_2_reg[14]  (.D(N239),
	.CLK(n25),
	.R(n55),
	.Q(result_2[14]));
   DFF \result_2_reg[13]  (.D(N238),
	.CLK(n20),
	.R(N0),
	.Q(result_2[13]));
   DFF \result_2_reg[12]  (.D(N237),
	.CLK(n22),
	.R(n54),
	.Q(result_2[12]));
   DFF \result_2_reg[11]  (.D(N236),
	.CLK(n57),
	.R(n55),
	.Q(result_2[11]));
   DFF \result_2_reg[10]  (.D(N235),
	.CLK(n60),
	.R(N0),
	.Q(result_2[10]));
   DFF \result_2_reg[9]  (.D(N234),
	.CLK(n58),
	.R(n54),
	.Q(result_2[9]));
   DFF \result_2_reg[8]  (.D(N233),
	.CLK(n29),
	.R(n55),
	.Q(result_2[8]));
   DFF \result_2_reg[7]  (.D(N232),
	.CLK(n18),
	.R(N0),
	.Q(result_2[7]));
   DFF \result_2_reg[6]  (.D(N231),
	.CLK(n27),
	.R(n54),
	.Q(result_2[6]));
   DFF \result_2_reg[5]  (.D(N230),
	.CLK(n37),
	.R(n55),
	.Q(result_2[5]));
   DFF \result_2_reg[4]  (.D(N229),
	.CLK(n65),
	.R(N0),
	.Q(result_2[4]));
   DFF \result_2_reg[3]  (.D(N228),
	.CLK(n36),
	.R(n54),
	.Q(result_2[3]));
   DFF \result_2_reg[2]  (.D(N227),
	.CLK(n19),
	.R(n55),
	.Q(result_2[2]));
   DFF \result_2_reg[1]  (.D(N226),
	.CLK(n41),
	.R(N0),
	.Q(result_2[1]));
   DFF \result_2_reg[0]  (.D(N225),
	.CLK(n26),
	.R(n54),
	.Q(result_2[0]));
   DFF \result_0_reg[15]  (.D(N80),
	.CLK(n24),
	.R(n55),
	.Q(result_0[15]));
   DFF \result_0_reg[14]  (.D(N79),
	.CLK(n42),
	.R(N0),
	.Q(result_0[14]));
   DFF \result_0_reg[13]  (.D(N78),
	.CLK(n50),
	.R(n54),
	.Q(result_0[13]));
   DFF \result_0_reg[12]  (.D(N77),
	.CLK(n63),
	.R(n55),
	.Q(result_0[12]));
   DFF \result_0_reg[11]  (.D(N76),
	.CLK(n59),
	.R(N0),
	.Q(result_0[11]));
   DFF \result_0_reg[10]  (.D(N75),
	.CLK(n35),
	.R(n54),
	.Q(result_0[10]));
   DFF \result_0_reg[9]  (.D(N74),
	.CLK(n31),
	.R(n55),
	.Q(result_0[9]));
   DFF \result_0_reg[8]  (.D(N73),
	.CLK(n30),
	.R(N0),
	.Q(result_0[8]));
   DFF \result_0_reg[7]  (.D(N72),
	.CLK(n49),
	.R(n54),
	.Q(result_0[7]));
   DFF \result_0_reg[6]  (.D(N71),
	.CLK(n51),
	.R(n55),
	.Q(result_0[6]));
   DFF \result_0_reg[5]  (.D(N70),
	.CLK(n46),
	.R(N0),
	.Q(result_0[5]));
   DFF \result_0_reg[4]  (.D(N69),
	.CLK(n64),
	.R(n54),
	.Q(result_0[4]));
   DFF \result_0_reg[3]  (.D(N68),
	.CLK(n48),
	.R(n55),
	.Q(result_0[3]));
   DFF \result_0_reg[2]  (.D(N67),
	.CLK(n56),
	.R(N0),
	.Q(result_0[2]));
   DFF \result_0_reg[1]  (.D(N66),
	.CLK(n62),
	.R(n54),
	.Q(result_0[1]));
   DFF \result_0_reg[0]  (.D(N65),
	.CLK(n33),
	.R(n55),
	.Q(result_0[0]));
   INVERTER U3 (.IN(clk),
	.OUT(n1));
   OAI21 \mult_21_3/FS_1/U6_1_0_3  (.OUT(\mult_21_3/FS_1/C[1][3][0] ),
	.C(n3329),
	.B(n3328),
	.A(n3327));
   OAI21 \mult_21_3/FS_1/U6_0_3_1  (.OUT(\mult_21_3/FS_1/C[1][3][1] ),
	.C(\mult_21_3/FS_1/G_n_int[0][3][0] ),
	.B(n3325),
	.A(n3324));
   XOR2 \mult_21_3/FS_1/U3_C_0_3_1  (.A(\mult_21_3/FS_1/PG_int[0][3][1] ),
	.B(\mult_21_3/FS_1/C[1][3][1] ),
	.OUT(N224));
   XOR2 \mult_21_3/FS_1/U3_C_0_3_0  (.A(\mult_21_3/FS_1/PG_int[0][3][0] ),
	.B(\mult_21_3/FS_1/C[1][3][0] ),
	.OUT(N223));
   NAND2 \mult_21_3/FS_1/U3_B_0_3_0  (.A(\mult_21_3/FS_1/G_n_int[0][3][0] ),
	.B(\mult_21_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3321));
   NAND2 \mult_21_3/FS_1/U2_0_3_0  (.A(\mult_21_3/A1[12] ),
	.B(\mult_21_3/A2[12] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_21_3/FS_1/U1_0_3_0  (.A(n3319),
	.B(n3320),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_21_3/FS_1/U6_0_2_3  (.OUT(\mult_21_3/FS_1/C[1][2][3] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][2] ),
	.B(n3318),
	.A(n3317));
   OAI21 \mult_21_3/FS_1/U5_0_2_3  (.OUT(\mult_21_3/FS_1/G[1][0][2] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][3] ),
	.B(n3316),
	.A(n3315));
   NAND2 \mult_21_3/FS_1/U4_0_2_3  (.A(\mult_21_3/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_21_3/FS_1/P[0][2][3] ),
	.OUT(n3328));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_3  (.A(\mult_21_3/FS_1/PG_int[0][2][3] ),
	.B(\mult_21_3/FS_1/C[1][2][3] ),
	.OUT(N222));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_3  (.A(\mult_21_3/FS_1/G_n_int[0][2][3] ),
	.B(\mult_21_3/FS_1/P[0][2][3] ),
	.OUT(n3314));
   NAND2 \mult_21_3/FS_1/U2_0_2_3  (.A(\mult_21_3/A1[11] ),
	.B(\mult_21_3/A2[11] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_3  (.A(n3312),
	.B(n3313),
	.OUT(\mult_21_3/FS_1/P[0][2][3] ));
   OAI21 \mult_21_3/FS_1/U6_0_2_2  (.OUT(\mult_21_3/FS_1/C[1][2][2] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][1] ),
	.B(n3311),
	.A(n3310));
   OAI21 \mult_21_3/FS_1/U5_0_2_2  (.OUT(\mult_21_3/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][2] ),
	.B(n3318),
	.A(n3309));
   NAND2 \mult_21_3/FS_1/U4_0_2_2  (.A(\mult_21_3/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_21_3/FS_1/P[0][2][2] ),
	.OUT(n3308));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_2  (.A(\mult_21_3/FS_1/PG_int[0][2][2] ),
	.B(\mult_21_3/FS_1/C[1][2][2] ),
	.OUT(N221));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_2  (.A(\mult_21_3/FS_1/G_n_int[0][2][2] ),
	.B(\mult_21_3/FS_1/P[0][2][2] ),
	.OUT(n3307));
   NAND2 \mult_21_3/FS_1/U2_0_2_2  (.A(\mult_21_3/A1[10] ),
	.B(\mult_21_3/A2[10] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_2  (.A(n3305),
	.B(n3306),
	.OUT(\mult_21_3/FS_1/P[0][2][2] ));
   OAI21 \mult_21_3/FS_1/U6_0_2_1  (.OUT(\mult_21_3/FS_1/C[1][2][1] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][0] ),
	.B(n3304),
	.A(n3327));
   OAI21 \mult_21_3/FS_1/U5_0_2_1  (.OUT(\mult_21_3/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_21_3/FS_1/G_n_int[0][2][1] ),
	.B(n3311),
	.A(\mult_21_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_3/FS_1/U4_0_2_1  (.A(\mult_21_3/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_21_3/FS_1/P[0][2][1] ),
	.OUT(n3303));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_1  (.A(\mult_21_3/FS_1/PG_int[0][2][1] ),
	.B(\mult_21_3/FS_1/C[1][2][1] ),
	.OUT(N220));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_1  (.A(\mult_21_3/FS_1/G_n_int[0][2][1] ),
	.B(\mult_21_3/FS_1/P[0][2][1] ),
	.OUT(n3302));
   NAND2 \mult_21_3/FS_1/U2_0_2_1  (.A(\mult_21_3/A1[9] ),
	.B(\mult_21_3/A2[9] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_1  (.A(n3300),
	.B(n3301),
	.OUT(\mult_21_3/FS_1/P[0][2][1] ));
   XOR2 \mult_21_3/FS_1/U3_C_0_2_0  (.A(\mult_21_3/FS_1/PG_int[0][2][0] ),
	.B(\mult_21_3/FS_1/C[1][2][0] ),
	.OUT(N219));
   NAND2 \mult_21_3/FS_1/U3_B_0_2_0  (.A(\mult_21_3/FS_1/G_n_int[0][2][0] ),
	.B(\mult_21_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3299));
   NAND2 \mult_21_3/FS_1/U2_0_2_0  (.A(\mult_21_3/A1[8] ),
	.B(\mult_21_3/A2[8] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_3/FS_1/U1_0_2_0  (.A(n3297),
	.B(n3298),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_21_3/FS_1/U3_B_0_1_3  (.A(\mult_21_3/FS_1/G_n_int[0][1][3] ),
	.B(\mult_21_3/FS_1/P[0][1][3] ),
	.OUT(n3296));
   NAND2 \mult_21_3/FS_1/U2_0_1_3  (.A(\mult_21_3/A1[7] ),
	.B(\mult_21_3/A2[7] ),
	.OUT(\mult_21_3/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_21_3/FS_1/U1_0_1_3  (.A(n3294),
	.B(n3295),
	.OUT(\mult_21_3/FS_1/P[0][1][3] ));
   INVERTER \mult_21_3/AN1_7  (.IN(matrix22[7]),
	.OUT(\mult_21_3/A_not[7] ));
   INVERTER \mult_21_3/AN1_6  (.IN(matrix22[6]),
	.OUT(\mult_21_3/A_notx [6]));
   INVERTER \mult_21_3/AN1_5  (.IN(matrix22[5]),
	.OUT(\mult_21_3/A_notx [5]));
   INVERTER \mult_21_3/AN1_4  (.IN(matrix22[4]),
	.OUT(\mult_21_3/A_notx [4]));
   INVERTER \mult_21_3/AN1_3  (.IN(matrix22[3]),
	.OUT(\mult_21_3/A_notx [3]));
   INVERTER \mult_21_3/AN1_2  (.IN(matrix22[2]),
	.OUT(\mult_21_3/A_notx [2]));
   INVERTER \mult_21_3/AN1_1  (.IN(matrix22[1]),
	.OUT(\mult_21_3/A_notx [1]));
   INVERTER \mult_21_3/AN1_0  (.IN(matrix22[0]),
	.OUT(\mult_21_3/A_notx [0]));
   INVERTER \mult_21_3/AN1_7_0  (.IN(vector_2[7]),
	.OUT(\mult_21_3/B_not[7] ));
   INVERTER \mult_21_3/AN1_6_0  (.IN(vector_2[6]),
	.OUT(\mult_21_3/B_notx [6]));
   INVERTER \mult_21_3/AN1_5_0  (.IN(vector_2[5]),
	.OUT(\mult_21_3/B_notx [5]));
   INVERTER \mult_21_3/AN1_4_0  (.IN(vector_2[4]),
	.OUT(\mult_21_3/B_notx [4]));
   INVERTER \mult_21_3/AN1_3_0  (.IN(vector_2[3]),
	.OUT(\mult_21_3/B_notx [3]));
   INVERTER \mult_21_3/AN1_2_0  (.IN(vector_2[2]),
	.OUT(\mult_21_3/B_notx [2]));
   INVERTER \mult_21_3/AN1_1_0  (.IN(vector_2[1]),
	.OUT(\mult_21_3/B_notx [1]));
   INVERTER \mult_21_3/AN1_0_0  (.IN(vector_2[0]),
	.OUT(\mult_21_3/B_notx [0]));
   NOR2 \mult_21_3/AN1_7_7  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[7][7] ));
   NOR2 \mult_21_3/AN3_7_6  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[7][6] ));
   NOR2 \mult_21_3/AN3_7_5  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[7][5] ));
   NOR2 \mult_21_3/AN3_7_4  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[7][4] ));
   NOR2 \mult_21_3/AN3_7_3  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[7][3] ));
   NOR2 \mult_21_3/AN3_7_2  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[7][2] ));
   NOR2 \mult_21_3/AN3_7_1  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[7][1] ));
   NOR2 \mult_21_3/AN3_7_0  (.A(\mult_21_3/A_not[7] ),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[7][0] ));
   NOR2 \mult_21_3/AN2_6_7  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[6][7] ));
   NOR2 \mult_21_3/AN1_6_6  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[6][6] ));
   NOR2 \mult_21_3/AN1_6_5  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[6][5] ));
   NOR2 \mult_21_3/AN1_6_4  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[6][4] ));
   NOR2 \mult_21_3/AN1_6_3  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[6][3] ));
   NOR2 \mult_21_3/AN1_6_2  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[6][2] ));
   NOR2 \mult_21_3/AN1_6_1  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[6][1] ));
   NOR2 \mult_21_3/AN1_6_0_0  (.A(\mult_21_3/A_notx [6]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[6][0] ));
   NOR2 \mult_21_3/AN2_5_7  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[5][7] ));
   NOR2 \mult_21_3/AN1_5_6  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[5][6] ));
   NOR2 \mult_21_3/AN1_5_5  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[5][5] ));
   NOR2 \mult_21_3/AN1_5_4  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[5][4] ));
   NOR2 \mult_21_3/AN1_5_3  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[5][3] ));
   NOR2 \mult_21_3/AN1_5_2  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[5][2] ));
   NOR2 \mult_21_3/AN1_5_1  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[5][1] ));
   NOR2 \mult_21_3/AN1_5_0_0  (.A(\mult_21_3/A_notx [5]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[5][0] ));
   NOR2 \mult_21_3/AN2_4_7  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[4][7] ));
   NOR2 \mult_21_3/AN1_4_6  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[4][6] ));
   NOR2 \mult_21_3/AN1_4_5  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[4][5] ));
   NOR2 \mult_21_3/AN1_4_4  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[4][4] ));
   NOR2 \mult_21_3/AN1_4_3  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[4][3] ));
   NOR2 \mult_21_3/AN1_4_2  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[4][2] ));
   NOR2 \mult_21_3/AN1_4_1  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[4][1] ));
   NOR2 \mult_21_3/AN1_4_0_0  (.A(\mult_21_3/A_notx [4]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[4][0] ));
   NOR2 \mult_21_3/AN2_3_7  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[3][7] ));
   NOR2 \mult_21_3/AN1_3_6  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[3][6] ));
   NOR2 \mult_21_3/AN1_3_5  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[3][5] ));
   NOR2 \mult_21_3/AN1_3_4  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[3][4] ));
   NOR2 \mult_21_3/AN1_3_3  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[3][3] ));
   NOR2 \mult_21_3/AN1_3_2  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[3][2] ));
   NOR2 \mult_21_3/AN1_3_1  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[3][1] ));
   NOR2 \mult_21_3/AN1_3_0_0  (.A(\mult_21_3/A_notx [3]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[3][0] ));
   NOR2 \mult_21_3/AN2_2_7  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[2][7] ));
   NOR2 \mult_21_3/AN1_2_6  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[2][6] ));
   NOR2 \mult_21_3/AN1_2_5  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[2][5] ));
   NOR2 \mult_21_3/AN1_2_4  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[2][4] ));
   NOR2 \mult_21_3/AN1_2_3  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[2][3] ));
   NOR2 \mult_21_3/AN1_2_2  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[2][2] ));
   NOR2 \mult_21_3/AN1_2_1  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[2][1] ));
   NOR2 \mult_21_3/AN1_2_0_0  (.A(\mult_21_3/A_notx [2]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[2][0] ));
   NOR2 \mult_21_3/AN2_1_7  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[1][7] ));
   NOR2 \mult_21_3/AN1_1_6  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[1][6] ));
   NOR2 \mult_21_3/AN1_1_5  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[1][5] ));
   NOR2 \mult_21_3/AN1_1_4  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[1][4] ));
   NOR2 \mult_21_3/AN1_1_3  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[1][3] ));
   NOR2 \mult_21_3/AN1_1_2  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[1][2] ));
   NOR2 \mult_21_3/AN1_1_1  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[1][1] ));
   NOR2 \mult_21_3/AN1_1_0_0  (.A(\mult_21_3/A_notx [1]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(\mult_21_3/ab[1][0] ));
   NOR2 \mult_21_3/AN2_0_7  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_not[7] ),
	.OUT(\mult_21_3/ab[0][7] ));
   NOR2 \mult_21_3/AN1_0_6  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [6]),
	.OUT(\mult_21_3/ab[0][6] ));
   NOR2 \mult_21_3/AN1_0_5  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [5]),
	.OUT(\mult_21_3/ab[0][5] ));
   NOR2 \mult_21_3/AN1_0_4  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [4]),
	.OUT(\mult_21_3/ab[0][4] ));
   NOR2 \mult_21_3/AN1_0_3  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [3]),
	.OUT(\mult_21_3/ab[0][3] ));
   NOR2 \mult_21_3/AN1_0_2  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [2]),
	.OUT(\mult_21_3/ab[0][2] ));
   NOR2 \mult_21_3/AN1_0_1  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [1]),
	.OUT(\mult_21_3/ab[0][1] ));
   NOR2 \mult_21_3/AN1_0_0_0  (.A(\mult_21_3/A_notx [0]),
	.B(\mult_21_3/B_notx [0]),
	.OUT(N209));
   OAI21 \mult_21_2/FS_1/U6_1_0_3  (.OUT(\mult_21_2/FS_1/C[1][3][0] ),
	.C(n3279),
	.B(n3278),
	.A(n3277));
   OAI21 \mult_21_2/FS_1/U6_0_3_1  (.OUT(\mult_21_2/FS_1/C[1][3][1] ),
	.C(\mult_21_2/FS_1/G_n_int[0][3][0] ),
	.B(n3275),
	.A(n3274));
   XOR2 \mult_21_2/FS_1/U3_C_0_3_1  (.A(\mult_21_2/FS_1/PG_int[0][3][1] ),
	.B(\mult_21_2/FS_1/C[1][3][1] ),
	.OUT(N192));
   XOR2 \mult_21_2/FS_1/U3_C_0_3_0  (.A(\mult_21_2/FS_1/PG_int[0][3][0] ),
	.B(\mult_21_2/FS_1/C[1][3][0] ),
	.OUT(N191));
   NAND2 \mult_21_2/FS_1/U3_B_0_3_0  (.A(\mult_21_2/FS_1/G_n_int[0][3][0] ),
	.B(\mult_21_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3271));
   NAND2 \mult_21_2/FS_1/U2_0_3_0  (.A(\mult_21_2/A1[12] ),
	.B(\mult_21_2/A2[12] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_21_2/FS_1/U1_0_3_0  (.A(n3269),
	.B(n3270),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_21_2/FS_1/U6_0_2_3  (.OUT(\mult_21_2/FS_1/C[1][2][3] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][2] ),
	.B(n3268),
	.A(n3267));
   OAI21 \mult_21_2/FS_1/U5_0_2_3  (.OUT(\mult_21_2/FS_1/G[1][0][2] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][3] ),
	.B(n3266),
	.A(n3265));
   NAND2 \mult_21_2/FS_1/U4_0_2_3  (.A(\mult_21_2/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_21_2/FS_1/P[0][2][3] ),
	.OUT(n3278));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_3  (.A(\mult_21_2/FS_1/PG_int[0][2][3] ),
	.B(\mult_21_2/FS_1/C[1][2][3] ),
	.OUT(N190));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_3  (.A(\mult_21_2/FS_1/G_n_int[0][2][3] ),
	.B(\mult_21_2/FS_1/P[0][2][3] ),
	.OUT(n3264));
   NAND2 \mult_21_2/FS_1/U2_0_2_3  (.A(\mult_21_2/A1[11] ),
	.B(\mult_21_2/A2[11] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_3  (.A(n3262),
	.B(n3263),
	.OUT(\mult_21_2/FS_1/P[0][2][3] ));
   OAI21 \mult_21_2/FS_1/U6_0_2_2  (.OUT(\mult_21_2/FS_1/C[1][2][2] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][1] ),
	.B(n3261),
	.A(n3260));
   OAI21 \mult_21_2/FS_1/U5_0_2_2  (.OUT(\mult_21_2/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][2] ),
	.B(n3268),
	.A(n3259));
   NAND2 \mult_21_2/FS_1/U4_0_2_2  (.A(\mult_21_2/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_21_2/FS_1/P[0][2][2] ),
	.OUT(n3258));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_2  (.A(\mult_21_2/FS_1/PG_int[0][2][2] ),
	.B(\mult_21_2/FS_1/C[1][2][2] ),
	.OUT(N189));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_2  (.A(\mult_21_2/FS_1/G_n_int[0][2][2] ),
	.B(\mult_21_2/FS_1/P[0][2][2] ),
	.OUT(n3257));
   NAND2 \mult_21_2/FS_1/U2_0_2_2  (.A(\mult_21_2/A1[10] ),
	.B(\mult_21_2/A2[10] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_2  (.A(n3255),
	.B(n3256),
	.OUT(\mult_21_2/FS_1/P[0][2][2] ));
   OAI21 \mult_21_2/FS_1/U6_0_2_1  (.OUT(\mult_21_2/FS_1/C[1][2][1] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][0] ),
	.B(n3254),
	.A(n3277));
   OAI21 \mult_21_2/FS_1/U5_0_2_1  (.OUT(\mult_21_2/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_21_2/FS_1/G_n_int[0][2][1] ),
	.B(n3261),
	.A(\mult_21_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_2/FS_1/U4_0_2_1  (.A(\mult_21_2/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_21_2/FS_1/P[0][2][1] ),
	.OUT(n3253));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_1  (.A(\mult_21_2/FS_1/PG_int[0][2][1] ),
	.B(\mult_21_2/FS_1/C[1][2][1] ),
	.OUT(N188));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_1  (.A(\mult_21_2/FS_1/G_n_int[0][2][1] ),
	.B(\mult_21_2/FS_1/P[0][2][1] ),
	.OUT(n3252));
   NAND2 \mult_21_2/FS_1/U2_0_2_1  (.A(\mult_21_2/A1[9] ),
	.B(\mult_21_2/A2[9] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_1  (.A(n3250),
	.B(n3251),
	.OUT(\mult_21_2/FS_1/P[0][2][1] ));
   XOR2 \mult_21_2/FS_1/U3_C_0_2_0  (.A(\mult_21_2/FS_1/PG_int[0][2][0] ),
	.B(\mult_21_2/FS_1/C[1][2][0] ),
	.OUT(N187));
   NAND2 \mult_21_2/FS_1/U3_B_0_2_0  (.A(\mult_21_2/FS_1/G_n_int[0][2][0] ),
	.B(\mult_21_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3249));
   NAND2 \mult_21_2/FS_1/U2_0_2_0  (.A(\mult_21_2/A1[8] ),
	.B(\mult_21_2/A2[8] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21_2/FS_1/U1_0_2_0  (.A(n3247),
	.B(n3248),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_21_2/FS_1/U3_B_0_1_3  (.A(\mult_21_2/FS_1/G_n_int[0][1][3] ),
	.B(\mult_21_2/FS_1/P[0][1][3] ),
	.OUT(n3246));
   NAND2 \mult_21_2/FS_1/U2_0_1_3  (.A(\mult_21_2/A1[7] ),
	.B(\mult_21_2/A2[7] ),
	.OUT(\mult_21_2/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_21_2/FS_1/U1_0_1_3  (.A(n3244),
	.B(n3245),
	.OUT(\mult_21_2/FS_1/P[0][1][3] ));
   INVERTER \mult_21_2/AN1_7  (.IN(matrix21[7]),
	.OUT(\mult_21_2/A_not[7] ));
   INVERTER \mult_21_2/AN1_6  (.IN(matrix21[6]),
	.OUT(\mult_21_2/A_notx [6]));
   INVERTER \mult_21_2/AN1_5  (.IN(matrix21[5]),
	.OUT(\mult_21_2/A_notx [5]));
   INVERTER \mult_21_2/AN1_4  (.IN(matrix21[4]),
	.OUT(\mult_21_2/A_notx [4]));
   INVERTER \mult_21_2/AN1_3  (.IN(matrix21[3]),
	.OUT(\mult_21_2/A_notx [3]));
   INVERTER \mult_21_2/AN1_2  (.IN(matrix21[2]),
	.OUT(\mult_21_2/A_notx [2]));
   INVERTER \mult_21_2/AN1_1  (.IN(matrix21[1]),
	.OUT(\mult_21_2/A_notx [1]));
   INVERTER \mult_21_2/AN1_0  (.IN(matrix21[0]),
	.OUT(\mult_21_2/A_notx [0]));
   INVERTER \mult_21_2/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_21_2/B_not[7] ));
   INVERTER \mult_21_2/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_21_2/B_notx [6]));
   INVERTER \mult_21_2/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_21_2/B_notx [5]));
   INVERTER \mult_21_2/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_21_2/B_notx [4]));
   INVERTER \mult_21_2/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_21_2/B_notx [3]));
   INVERTER \mult_21_2/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_21_2/B_notx [2]));
   INVERTER \mult_21_2/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_21_2/B_notx [1]));
   INVERTER \mult_21_2/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_21_2/B_notx [0]));
   NOR2 \mult_21_2/AN1_7_7  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[7][7] ));
   NOR2 \mult_21_2/AN3_7_6  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[7][6] ));
   NOR2 \mult_21_2/AN3_7_5  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[7][5] ));
   NOR2 \mult_21_2/AN3_7_4  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[7][4] ));
   NOR2 \mult_21_2/AN3_7_3  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[7][3] ));
   NOR2 \mult_21_2/AN3_7_2  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[7][2] ));
   NOR2 \mult_21_2/AN3_7_1  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[7][1] ));
   NOR2 \mult_21_2/AN3_7_0  (.A(\mult_21_2/A_not[7] ),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[7][0] ));
   NOR2 \mult_21_2/AN2_6_7  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[6][7] ));
   NOR2 \mult_21_2/AN1_6_6  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[6][6] ));
   NOR2 \mult_21_2/AN1_6_5  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[6][5] ));
   NOR2 \mult_21_2/AN1_6_4  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[6][4] ));
   NOR2 \mult_21_2/AN1_6_3  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[6][3] ));
   NOR2 \mult_21_2/AN1_6_2  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[6][2] ));
   NOR2 \mult_21_2/AN1_6_1  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[6][1] ));
   NOR2 \mult_21_2/AN1_6_0_0  (.A(\mult_21_2/A_notx [6]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[6][0] ));
   NOR2 \mult_21_2/AN2_5_7  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[5][7] ));
   NOR2 \mult_21_2/AN1_5_6  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[5][6] ));
   NOR2 \mult_21_2/AN1_5_5  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[5][5] ));
   NOR2 \mult_21_2/AN1_5_4  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[5][4] ));
   NOR2 \mult_21_2/AN1_5_3  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[5][3] ));
   NOR2 \mult_21_2/AN1_5_2  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[5][2] ));
   NOR2 \mult_21_2/AN1_5_1  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[5][1] ));
   NOR2 \mult_21_2/AN1_5_0_0  (.A(\mult_21_2/A_notx [5]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[5][0] ));
   NOR2 \mult_21_2/AN2_4_7  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[4][7] ));
   NOR2 \mult_21_2/AN1_4_6  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[4][6] ));
   NOR2 \mult_21_2/AN1_4_5  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[4][5] ));
   NOR2 \mult_21_2/AN1_4_4  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[4][4] ));
   NOR2 \mult_21_2/AN1_4_3  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[4][3] ));
   NOR2 \mult_21_2/AN1_4_2  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[4][2] ));
   NOR2 \mult_21_2/AN1_4_1  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[4][1] ));
   NOR2 \mult_21_2/AN1_4_0_0  (.A(\mult_21_2/A_notx [4]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[4][0] ));
   NOR2 \mult_21_2/AN2_3_7  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[3][7] ));
   NOR2 \mult_21_2/AN1_3_6  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[3][6] ));
   NOR2 \mult_21_2/AN1_3_5  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[3][5] ));
   NOR2 \mult_21_2/AN1_3_4  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[3][4] ));
   NOR2 \mult_21_2/AN1_3_3  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[3][3] ));
   NOR2 \mult_21_2/AN1_3_2  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[3][2] ));
   NOR2 \mult_21_2/AN1_3_1  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[3][1] ));
   NOR2 \mult_21_2/AN1_3_0_0  (.A(\mult_21_2/A_notx [3]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[3][0] ));
   NOR2 \mult_21_2/AN2_2_7  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[2][7] ));
   NOR2 \mult_21_2/AN1_2_6  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[2][6] ));
   NOR2 \mult_21_2/AN1_2_5  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[2][5] ));
   NOR2 \mult_21_2/AN1_2_4  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[2][4] ));
   NOR2 \mult_21_2/AN1_2_3  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[2][3] ));
   NOR2 \mult_21_2/AN1_2_2  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[2][2] ));
   NOR2 \mult_21_2/AN1_2_1  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[2][1] ));
   NOR2 \mult_21_2/AN1_2_0_0  (.A(\mult_21_2/A_notx [2]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[2][0] ));
   NOR2 \mult_21_2/AN2_1_7  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[1][7] ));
   NOR2 \mult_21_2/AN1_1_6  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[1][6] ));
   NOR2 \mult_21_2/AN1_1_5  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[1][5] ));
   NOR2 \mult_21_2/AN1_1_4  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[1][4] ));
   NOR2 \mult_21_2/AN1_1_3  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[1][3] ));
   NOR2 \mult_21_2/AN1_1_2  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[1][2] ));
   NOR2 \mult_21_2/AN1_1_1  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[1][1] ));
   NOR2 \mult_21_2/AN1_1_0_0  (.A(\mult_21_2/A_notx [1]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(\mult_21_2/ab[1][0] ));
   NOR2 \mult_21_2/AN2_0_7  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_not[7] ),
	.OUT(\mult_21_2/ab[0][7] ));
   NOR2 \mult_21_2/AN1_0_6  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [6]),
	.OUT(\mult_21_2/ab[0][6] ));
   NOR2 \mult_21_2/AN1_0_5  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [5]),
	.OUT(\mult_21_2/ab[0][5] ));
   NOR2 \mult_21_2/AN1_0_4  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [4]),
	.OUT(\mult_21_2/ab[0][4] ));
   NOR2 \mult_21_2/AN1_0_3  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [3]),
	.OUT(\mult_21_2/ab[0][3] ));
   NOR2 \mult_21_2/AN1_0_2  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [2]),
	.OUT(\mult_21_2/ab[0][2] ));
   NOR2 \mult_21_2/AN1_0_1  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [1]),
	.OUT(\mult_21_2/ab[0][1] ));
   NOR2 \mult_21_2/AN1_0_0_0  (.A(\mult_21_2/A_notx [0]),
	.B(\mult_21_2/B_notx [0]),
	.OUT(N177));
   OAI21 \mult_21/FS_1/U6_1_0_3  (.OUT(\mult_21/FS_1/C[1][3][0] ),
	.C(n3229),
	.B(n3228),
	.A(n3227));
   OAI21 \mult_21/FS_1/U6_0_3_1  (.OUT(\mult_21/FS_1/C[1][3][1] ),
	.C(\mult_21/FS_1/G_n_int[0][3][0] ),
	.B(n3225),
	.A(n3224));
   XOR2 \mult_21/FS_1/U3_C_0_3_1  (.A(\mult_21/FS_1/PG_int[0][3][1] ),
	.B(\mult_21/FS_1/C[1][3][1] ),
	.OUT(N176));
   XOR2 \mult_21/FS_1/U3_C_0_3_0  (.A(\mult_21/FS_1/PG_int[0][3][0] ),
	.B(\mult_21/FS_1/C[1][3][0] ),
	.OUT(N175));
   NAND2 \mult_21/FS_1/U3_B_0_3_0  (.A(\mult_21/FS_1/G_n_int[0][3][0] ),
	.B(\mult_21/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3221));
   NAND2 \mult_21/FS_1/U2_0_3_0  (.A(\mult_21/A1[12] ),
	.B(\mult_21/A2[12] ),
	.OUT(\mult_21/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_21/FS_1/U1_0_3_0  (.A(n3219),
	.B(n3220),
	.OUT(\mult_21/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_21/FS_1/U6_0_2_3  (.OUT(\mult_21/FS_1/C[1][2][3] ),
	.C(\mult_21/FS_1/G_n_int[0][2][2] ),
	.B(n3218),
	.A(n3217));
   OAI21 \mult_21/FS_1/U5_0_2_3  (.OUT(\mult_21/FS_1/G[1][0][2] ),
	.C(\mult_21/FS_1/G_n_int[0][2][3] ),
	.B(n3216),
	.A(n3215));
   NAND2 \mult_21/FS_1/U4_0_2_3  (.A(\mult_21/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_21/FS_1/P[0][2][3] ),
	.OUT(n3228));
   XOR2 \mult_21/FS_1/U3_C_0_2_3  (.A(\mult_21/FS_1/PG_int[0][2][3] ),
	.B(\mult_21/FS_1/C[1][2][3] ),
	.OUT(N174));
   NAND2 \mult_21/FS_1/U3_B_0_2_3  (.A(\mult_21/FS_1/G_n_int[0][2][3] ),
	.B(\mult_21/FS_1/P[0][2][3] ),
	.OUT(n3214));
   NAND2 \mult_21/FS_1/U2_0_2_3  (.A(\mult_21/A1[11] ),
	.B(\mult_21/A2[11] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_21/FS_1/U1_0_2_3  (.A(n3212),
	.B(n3213),
	.OUT(\mult_21/FS_1/P[0][2][3] ));
   OAI21 \mult_21/FS_1/U6_0_2_2  (.OUT(\mult_21/FS_1/C[1][2][2] ),
	.C(\mult_21/FS_1/G_n_int[0][2][1] ),
	.B(n3211),
	.A(n3210));
   OAI21 \mult_21/FS_1/U5_0_2_2  (.OUT(\mult_21/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_21/FS_1/G_n_int[0][2][2] ),
	.B(n3218),
	.A(n3209));
   NAND2 \mult_21/FS_1/U4_0_2_2  (.A(\mult_21/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_21/FS_1/P[0][2][2] ),
	.OUT(n3208));
   XOR2 \mult_21/FS_1/U3_C_0_2_2  (.A(\mult_21/FS_1/PG_int[0][2][2] ),
	.B(\mult_21/FS_1/C[1][2][2] ),
	.OUT(N173));
   NAND2 \mult_21/FS_1/U3_B_0_2_2  (.A(\mult_21/FS_1/G_n_int[0][2][2] ),
	.B(\mult_21/FS_1/P[0][2][2] ),
	.OUT(n3207));
   NAND2 \mult_21/FS_1/U2_0_2_2  (.A(\mult_21/A1[10] ),
	.B(\mult_21/A2[10] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_21/FS_1/U1_0_2_2  (.A(n3205),
	.B(n3206),
	.OUT(\mult_21/FS_1/P[0][2][2] ));
   OAI21 \mult_21/FS_1/U6_0_2_1  (.OUT(\mult_21/FS_1/C[1][2][1] ),
	.C(\mult_21/FS_1/G_n_int[0][2][0] ),
	.B(n3204),
	.A(n3227));
   OAI21 \mult_21/FS_1/U5_0_2_1  (.OUT(\mult_21/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_21/FS_1/G_n_int[0][2][1] ),
	.B(n3211),
	.A(\mult_21/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21/FS_1/U4_0_2_1  (.A(\mult_21/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_21/FS_1/P[0][2][1] ),
	.OUT(n3203));
   XOR2 \mult_21/FS_1/U3_C_0_2_1  (.A(\mult_21/FS_1/PG_int[0][2][1] ),
	.B(\mult_21/FS_1/C[1][2][1] ),
	.OUT(N172));
   NAND2 \mult_21/FS_1/U3_B_0_2_1  (.A(\mult_21/FS_1/G_n_int[0][2][1] ),
	.B(\mult_21/FS_1/P[0][2][1] ),
	.OUT(n3202));
   NAND2 \mult_21/FS_1/U2_0_2_1  (.A(\mult_21/A1[9] ),
	.B(\mult_21/A2[9] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_21/FS_1/U1_0_2_1  (.A(n3200),
	.B(n3201),
	.OUT(\mult_21/FS_1/P[0][2][1] ));
   XOR2 \mult_21/FS_1/U3_C_0_2_0  (.A(\mult_21/FS_1/PG_int[0][2][0] ),
	.B(\mult_21/FS_1/C[1][2][0] ),
	.OUT(N171));
   NAND2 \mult_21/FS_1/U3_B_0_2_0  (.A(\mult_21/FS_1/G_n_int[0][2][0] ),
	.B(\mult_21/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3199));
   NAND2 \mult_21/FS_1/U2_0_2_0  (.A(\mult_21/A1[8] ),
	.B(\mult_21/A2[8] ),
	.OUT(\mult_21/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_21/FS_1/U1_0_2_0  (.A(n3197),
	.B(n3198),
	.OUT(\mult_21/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_21/FS_1/U3_B_0_1_3  (.A(\mult_21/FS_1/G_n_int[0][1][3] ),
	.B(\mult_21/FS_1/P[0][1][3] ),
	.OUT(n3196));
   NAND2 \mult_21/FS_1/U2_0_1_3  (.A(\mult_21/A1[7] ),
	.B(\mult_21/A2[7] ),
	.OUT(\mult_21/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_21/FS_1/U1_0_1_3  (.A(n3194),
	.B(n3195),
	.OUT(\mult_21/FS_1/P[0][1][3] ));
   INVERTER \mult_21/AN1_7  (.IN(matrix20[7]),
	.OUT(\mult_21/A_not[7] ));
   INVERTER \mult_21/AN1_6  (.IN(matrix20[6]),
	.OUT(\mult_21/A_notx [6]));
   INVERTER \mult_21/AN1_5  (.IN(matrix20[5]),
	.OUT(\mult_21/A_notx [5]));
   INVERTER \mult_21/AN1_4  (.IN(matrix20[4]),
	.OUT(\mult_21/A_notx [4]));
   INVERTER \mult_21/AN1_3  (.IN(matrix20[3]),
	.OUT(\mult_21/A_notx [3]));
   INVERTER \mult_21/AN1_2  (.IN(matrix20[2]),
	.OUT(\mult_21/A_notx [2]));
   INVERTER \mult_21/AN1_1  (.IN(matrix20[1]),
	.OUT(\mult_21/A_notx [1]));
   INVERTER \mult_21/AN1_0  (.IN(matrix20[0]),
	.OUT(\mult_21/A_notx [0]));
   INVERTER \mult_21/AN1_7_0  (.IN(vector_0[7]),
	.OUT(\mult_21/B_not[7] ));
   INVERTER \mult_21/AN1_6_0  (.IN(vector_0[6]),
	.OUT(\mult_21/B_notx [6]));
   INVERTER \mult_21/AN1_5_0  (.IN(vector_0[5]),
	.OUT(\mult_21/B_notx [5]));
   INVERTER \mult_21/AN1_4_0  (.IN(vector_0[4]),
	.OUT(\mult_21/B_notx [4]));
   INVERTER \mult_21/AN1_3_0  (.IN(vector_0[3]),
	.OUT(\mult_21/B_notx [3]));
   INVERTER \mult_21/AN1_2_0  (.IN(vector_0[2]),
	.OUT(\mult_21/B_notx [2]));
   INVERTER \mult_21/AN1_1_0  (.IN(vector_0[1]),
	.OUT(\mult_21/B_notx [1]));
   INVERTER \mult_21/AN1_0_0  (.IN(vector_0[0]),
	.OUT(\mult_21/B_notx [0]));
   NOR2 \mult_21/AN1_7_7  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[7][7] ));
   NOR2 \mult_21/AN3_7_6  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[7][6] ));
   NOR2 \mult_21/AN3_7_5  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[7][5] ));
   NOR2 \mult_21/AN3_7_4  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[7][4] ));
   NOR2 \mult_21/AN3_7_3  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[7][3] ));
   NOR2 \mult_21/AN3_7_2  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[7][2] ));
   NOR2 \mult_21/AN3_7_1  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[7][1] ));
   NOR2 \mult_21/AN3_7_0  (.A(\mult_21/A_not[7] ),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[7][0] ));
   NOR2 \mult_21/AN2_6_7  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[6][7] ));
   NOR2 \mult_21/AN1_6_6  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[6][6] ));
   NOR2 \mult_21/AN1_6_5  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[6][5] ));
   NOR2 \mult_21/AN1_6_4  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[6][4] ));
   NOR2 \mult_21/AN1_6_3  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[6][3] ));
   NOR2 \mult_21/AN1_6_2  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[6][2] ));
   NOR2 \mult_21/AN1_6_1  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[6][1] ));
   NOR2 \mult_21/AN1_6_0_0  (.A(\mult_21/A_notx [6]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[6][0] ));
   NOR2 \mult_21/AN2_5_7  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[5][7] ));
   NOR2 \mult_21/AN1_5_6  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[5][6] ));
   NOR2 \mult_21/AN1_5_5  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[5][5] ));
   NOR2 \mult_21/AN1_5_4  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[5][4] ));
   NOR2 \mult_21/AN1_5_3  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[5][3] ));
   NOR2 \mult_21/AN1_5_2  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[5][2] ));
   NOR2 \mult_21/AN1_5_1  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[5][1] ));
   NOR2 \mult_21/AN1_5_0_0  (.A(\mult_21/A_notx [5]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[5][0] ));
   NOR2 \mult_21/AN2_4_7  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[4][7] ));
   NOR2 \mult_21/AN1_4_6  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[4][6] ));
   NOR2 \mult_21/AN1_4_5  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[4][5] ));
   NOR2 \mult_21/AN1_4_4  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[4][4] ));
   NOR2 \mult_21/AN1_4_3  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[4][3] ));
   NOR2 \mult_21/AN1_4_2  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[4][2] ));
   NOR2 \mult_21/AN1_4_1  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[4][1] ));
   NOR2 \mult_21/AN1_4_0_0  (.A(\mult_21/A_notx [4]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[4][0] ));
   NOR2 \mult_21/AN2_3_7  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[3][7] ));
   NOR2 \mult_21/AN1_3_6  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[3][6] ));
   NOR2 \mult_21/AN1_3_5  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[3][5] ));
   NOR2 \mult_21/AN1_3_4  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[3][4] ));
   NOR2 \mult_21/AN1_3_3  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[3][3] ));
   NOR2 \mult_21/AN1_3_2  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[3][2] ));
   NOR2 \mult_21/AN1_3_1  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[3][1] ));
   NOR2 \mult_21/AN1_3_0_0  (.A(\mult_21/A_notx [3]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[3][0] ));
   NOR2 \mult_21/AN2_2_7  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[2][7] ));
   NOR2 \mult_21/AN1_2_6  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[2][6] ));
   NOR2 \mult_21/AN1_2_5  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[2][5] ));
   NOR2 \mult_21/AN1_2_4  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[2][4] ));
   NOR2 \mult_21/AN1_2_3  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[2][3] ));
   NOR2 \mult_21/AN1_2_2  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[2][2] ));
   NOR2 \mult_21/AN1_2_1  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[2][1] ));
   NOR2 \mult_21/AN1_2_0_0  (.A(\mult_21/A_notx [2]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[2][0] ));
   NOR2 \mult_21/AN2_1_7  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[1][7] ));
   NOR2 \mult_21/AN1_1_6  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[1][6] ));
   NOR2 \mult_21/AN1_1_5  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[1][5] ));
   NOR2 \mult_21/AN1_1_4  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[1][4] ));
   NOR2 \mult_21/AN1_1_3  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[1][3] ));
   NOR2 \mult_21/AN1_1_2  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[1][2] ));
   NOR2 \mult_21/AN1_1_1  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[1][1] ));
   NOR2 \mult_21/AN1_1_0_0  (.A(\mult_21/A_notx [1]),
	.B(\mult_21/B_notx [0]),
	.OUT(\mult_21/ab[1][0] ));
   NOR2 \mult_21/AN2_0_7  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_not[7] ),
	.OUT(\mult_21/ab[0][7] ));
   NOR2 \mult_21/AN1_0_6  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [6]),
	.OUT(\mult_21/ab[0][6] ));
   NOR2 \mult_21/AN1_0_5  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [5]),
	.OUT(\mult_21/ab[0][5] ));
   NOR2 \mult_21/AN1_0_4  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [4]),
	.OUT(\mult_21/ab[0][4] ));
   NOR2 \mult_21/AN1_0_3  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [3]),
	.OUT(\mult_21/ab[0][3] ));
   NOR2 \mult_21/AN1_0_2  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [2]),
	.OUT(\mult_21/ab[0][2] ));
   NOR2 \mult_21/AN1_0_1  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [1]),
	.OUT(\mult_21/ab[0][1] ));
   NOR2 \mult_21/AN1_0_0_0  (.A(\mult_21/A_notx [0]),
	.B(\mult_21/B_notx [0]),
	.OUT(N161));
   OAI21 \mult_20_3/FS_1/U6_1_0_3  (.OUT(\mult_20_3/FS_1/C[1][3][0] ),
	.C(n3179),
	.B(n3178),
	.A(n3177));
   OAI21 \mult_20_3/FS_1/U6_0_3_1  (.OUT(\mult_20_3/FS_1/C[1][3][1] ),
	.C(\mult_20_3/FS_1/G_n_int[0][3][0] ),
	.B(n3175),
	.A(n3174));
   XOR2 \mult_20_3/FS_1/U3_C_0_3_1  (.A(\mult_20_3/FS_1/PG_int[0][3][1] ),
	.B(\mult_20_3/FS_1/C[1][3][1] ),
	.OUT(N144));
   XOR2 \mult_20_3/FS_1/U3_C_0_3_0  (.A(\mult_20_3/FS_1/PG_int[0][3][0] ),
	.B(\mult_20_3/FS_1/C[1][3][0] ),
	.OUT(N143));
   NAND2 \mult_20_3/FS_1/U3_B_0_3_0  (.A(\mult_20_3/FS_1/G_n_int[0][3][0] ),
	.B(\mult_20_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3171));
   NAND2 \mult_20_3/FS_1/U2_0_3_0  (.A(\mult_20_3/A1[12] ),
	.B(\mult_20_3/A2[12] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_20_3/FS_1/U1_0_3_0  (.A(n3169),
	.B(n3170),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_20_3/FS_1/U6_0_2_3  (.OUT(\mult_20_3/FS_1/C[1][2][3] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][2] ),
	.B(n3168),
	.A(n3167));
   OAI21 \mult_20_3/FS_1/U5_0_2_3  (.OUT(\mult_20_3/FS_1/G[1][0][2] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][3] ),
	.B(n3166),
	.A(n3165));
   NAND2 \mult_20_3/FS_1/U4_0_2_3  (.A(\mult_20_3/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_20_3/FS_1/P[0][2][3] ),
	.OUT(n3178));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_3  (.A(\mult_20_3/FS_1/PG_int[0][2][3] ),
	.B(\mult_20_3/FS_1/C[1][2][3] ),
	.OUT(N142));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_3  (.A(\mult_20_3/FS_1/G_n_int[0][2][3] ),
	.B(\mult_20_3/FS_1/P[0][2][3] ),
	.OUT(n3164));
   NAND2 \mult_20_3/FS_1/U2_0_2_3  (.A(\mult_20_3/A1[11] ),
	.B(\mult_20_3/A2[11] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_3  (.A(n3162),
	.B(n3163),
	.OUT(\mult_20_3/FS_1/P[0][2][3] ));
   OAI21 \mult_20_3/FS_1/U6_0_2_2  (.OUT(\mult_20_3/FS_1/C[1][2][2] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][1] ),
	.B(n3161),
	.A(n3160));
   OAI21 \mult_20_3/FS_1/U5_0_2_2  (.OUT(\mult_20_3/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][2] ),
	.B(n3168),
	.A(n3159));
   NAND2 \mult_20_3/FS_1/U4_0_2_2  (.A(\mult_20_3/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_20_3/FS_1/P[0][2][2] ),
	.OUT(n3158));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_2  (.A(\mult_20_3/FS_1/PG_int[0][2][2] ),
	.B(\mult_20_3/FS_1/C[1][2][2] ),
	.OUT(N141));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_2  (.A(\mult_20_3/FS_1/G_n_int[0][2][2] ),
	.B(\mult_20_3/FS_1/P[0][2][2] ),
	.OUT(n3157));
   NAND2 \mult_20_3/FS_1/U2_0_2_2  (.A(\mult_20_3/A1[10] ),
	.B(\mult_20_3/A2[10] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_2  (.A(n3155),
	.B(n3156),
	.OUT(\mult_20_3/FS_1/P[0][2][2] ));
   OAI21 \mult_20_3/FS_1/U6_0_2_1  (.OUT(\mult_20_3/FS_1/C[1][2][1] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][0] ),
	.B(n3154),
	.A(n3177));
   OAI21 \mult_20_3/FS_1/U5_0_2_1  (.OUT(\mult_20_3/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_20_3/FS_1/G_n_int[0][2][1] ),
	.B(n3161),
	.A(\mult_20_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_3/FS_1/U4_0_2_1  (.A(\mult_20_3/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_20_3/FS_1/P[0][2][1] ),
	.OUT(n3153));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_1  (.A(\mult_20_3/FS_1/PG_int[0][2][1] ),
	.B(\mult_20_3/FS_1/C[1][2][1] ),
	.OUT(N140));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_1  (.A(\mult_20_3/FS_1/G_n_int[0][2][1] ),
	.B(\mult_20_3/FS_1/P[0][2][1] ),
	.OUT(n3152));
   NAND2 \mult_20_3/FS_1/U2_0_2_1  (.A(\mult_20_3/A1[9] ),
	.B(\mult_20_3/A2[9] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_1  (.A(n3150),
	.B(n3151),
	.OUT(\mult_20_3/FS_1/P[0][2][1] ));
   XOR2 \mult_20_3/FS_1/U3_C_0_2_0  (.A(\mult_20_3/FS_1/PG_int[0][2][0] ),
	.B(\mult_20_3/FS_1/C[1][2][0] ),
	.OUT(N139));
   NAND2 \mult_20_3/FS_1/U3_B_0_2_0  (.A(\mult_20_3/FS_1/G_n_int[0][2][0] ),
	.B(\mult_20_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3149));
   NAND2 \mult_20_3/FS_1/U2_0_2_0  (.A(\mult_20_3/A1[8] ),
	.B(\mult_20_3/A2[8] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_3/FS_1/U1_0_2_0  (.A(n3147),
	.B(n3148),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_20_3/FS_1/U3_B_0_1_3  (.A(\mult_20_3/FS_1/G_n_int[0][1][3] ),
	.B(\mult_20_3/FS_1/P[0][1][3] ),
	.OUT(n3146));
   NAND2 \mult_20_3/FS_1/U2_0_1_3  (.A(\mult_20_3/A1[7] ),
	.B(\mult_20_3/A2[7] ),
	.OUT(\mult_20_3/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_20_3/FS_1/U1_0_1_3  (.A(n3144),
	.B(n3145),
	.OUT(\mult_20_3/FS_1/P[0][1][3] ));
   INVERTER \mult_20_3/AN1_7  (.IN(matrix12[7]),
	.OUT(\mult_20_3/A_not[7] ));
   INVERTER \mult_20_3/AN1_6  (.IN(matrix12[6]),
	.OUT(\mult_20_3/A_notx [6]));
   INVERTER \mult_20_3/AN1_5  (.IN(matrix12[5]),
	.OUT(\mult_20_3/A_notx [5]));
   INVERTER \mult_20_3/AN1_4  (.IN(matrix12[4]),
	.OUT(\mult_20_3/A_notx [4]));
   INVERTER \mult_20_3/AN1_3  (.IN(matrix12[3]),
	.OUT(\mult_20_3/A_notx [3]));
   INVERTER \mult_20_3/AN1_2  (.IN(matrix12[2]),
	.OUT(\mult_20_3/A_notx [2]));
   INVERTER \mult_20_3/AN1_1  (.IN(matrix12[1]),
	.OUT(\mult_20_3/A_notx [1]));
   INVERTER \mult_20_3/AN1_0  (.IN(matrix12[0]),
	.OUT(\mult_20_3/A_notx [0]));
   INVERTER \mult_20_3/AN1_7_0  (.IN(vector_2[7]),
	.OUT(\mult_20_3/B_not[7] ));
   INVERTER \mult_20_3/AN1_6_0  (.IN(vector_2[6]),
	.OUT(\mult_20_3/B_notx [6]));
   INVERTER \mult_20_3/AN1_5_0  (.IN(vector_2[5]),
	.OUT(\mult_20_3/B_notx [5]));
   INVERTER \mult_20_3/AN1_4_0  (.IN(vector_2[4]),
	.OUT(\mult_20_3/B_notx [4]));
   INVERTER \mult_20_3/AN1_3_0  (.IN(vector_2[3]),
	.OUT(\mult_20_3/B_notx [3]));
   INVERTER \mult_20_3/AN1_2_0  (.IN(vector_2[2]),
	.OUT(\mult_20_3/B_notx [2]));
   INVERTER \mult_20_3/AN1_1_0  (.IN(vector_2[1]),
	.OUT(\mult_20_3/B_notx [1]));
   INVERTER \mult_20_3/AN1_0_0  (.IN(vector_2[0]),
	.OUT(\mult_20_3/B_notx [0]));
   NOR2 \mult_20_3/AN1_7_7  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[7][7] ));
   NOR2 \mult_20_3/AN3_7_6  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[7][6] ));
   NOR2 \mult_20_3/AN3_7_5  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[7][5] ));
   NOR2 \mult_20_3/AN3_7_4  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[7][4] ));
   NOR2 \mult_20_3/AN3_7_3  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[7][3] ));
   NOR2 \mult_20_3/AN3_7_2  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[7][2] ));
   NOR2 \mult_20_3/AN3_7_1  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[7][1] ));
   NOR2 \mult_20_3/AN3_7_0  (.A(\mult_20_3/A_not[7] ),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[7][0] ));
   NOR2 \mult_20_3/AN2_6_7  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[6][7] ));
   NOR2 \mult_20_3/AN1_6_6  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[6][6] ));
   NOR2 \mult_20_3/AN1_6_5  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[6][5] ));
   NOR2 \mult_20_3/AN1_6_4  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[6][4] ));
   NOR2 \mult_20_3/AN1_6_3  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[6][3] ));
   NOR2 \mult_20_3/AN1_6_2  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[6][2] ));
   NOR2 \mult_20_3/AN1_6_1  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[6][1] ));
   NOR2 \mult_20_3/AN1_6_0_0  (.A(\mult_20_3/A_notx [6]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[6][0] ));
   NOR2 \mult_20_3/AN2_5_7  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[5][7] ));
   NOR2 \mult_20_3/AN1_5_6  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[5][6] ));
   NOR2 \mult_20_3/AN1_5_5  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[5][5] ));
   NOR2 \mult_20_3/AN1_5_4  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[5][4] ));
   NOR2 \mult_20_3/AN1_5_3  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[5][3] ));
   NOR2 \mult_20_3/AN1_5_2  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[5][2] ));
   NOR2 \mult_20_3/AN1_5_1  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[5][1] ));
   NOR2 \mult_20_3/AN1_5_0_0  (.A(\mult_20_3/A_notx [5]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[5][0] ));
   NOR2 \mult_20_3/AN2_4_7  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[4][7] ));
   NOR2 \mult_20_3/AN1_4_6  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[4][6] ));
   NOR2 \mult_20_3/AN1_4_5  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[4][5] ));
   NOR2 \mult_20_3/AN1_4_4  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[4][4] ));
   NOR2 \mult_20_3/AN1_4_3  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[4][3] ));
   NOR2 \mult_20_3/AN1_4_2  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[4][2] ));
   NOR2 \mult_20_3/AN1_4_1  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[4][1] ));
   NOR2 \mult_20_3/AN1_4_0_0  (.A(\mult_20_3/A_notx [4]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[4][0] ));
   NOR2 \mult_20_3/AN2_3_7  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[3][7] ));
   NOR2 \mult_20_3/AN1_3_6  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[3][6] ));
   NOR2 \mult_20_3/AN1_3_5  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[3][5] ));
   NOR2 \mult_20_3/AN1_3_4  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[3][4] ));
   NOR2 \mult_20_3/AN1_3_3  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[3][3] ));
   NOR2 \mult_20_3/AN1_3_2  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[3][2] ));
   NOR2 \mult_20_3/AN1_3_1  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[3][1] ));
   NOR2 \mult_20_3/AN1_3_0_0  (.A(\mult_20_3/A_notx [3]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[3][0] ));
   NOR2 \mult_20_3/AN2_2_7  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[2][7] ));
   NOR2 \mult_20_3/AN1_2_6  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[2][6] ));
   NOR2 \mult_20_3/AN1_2_5  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[2][5] ));
   NOR2 \mult_20_3/AN1_2_4  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[2][4] ));
   NOR2 \mult_20_3/AN1_2_3  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[2][3] ));
   NOR2 \mult_20_3/AN1_2_2  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[2][2] ));
   NOR2 \mult_20_3/AN1_2_1  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[2][1] ));
   NOR2 \mult_20_3/AN1_2_0_0  (.A(\mult_20_3/A_notx [2]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[2][0] ));
   NOR2 \mult_20_3/AN2_1_7  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[1][7] ));
   NOR2 \mult_20_3/AN1_1_6  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[1][6] ));
   NOR2 \mult_20_3/AN1_1_5  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[1][5] ));
   NOR2 \mult_20_3/AN1_1_4  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[1][4] ));
   NOR2 \mult_20_3/AN1_1_3  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[1][3] ));
   NOR2 \mult_20_3/AN1_1_2  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[1][2] ));
   NOR2 \mult_20_3/AN1_1_1  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[1][1] ));
   NOR2 \mult_20_3/AN1_1_0_0  (.A(\mult_20_3/A_notx [1]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(\mult_20_3/ab[1][0] ));
   NOR2 \mult_20_3/AN2_0_7  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_not[7] ),
	.OUT(\mult_20_3/ab[0][7] ));
   NOR2 \mult_20_3/AN1_0_6  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [6]),
	.OUT(\mult_20_3/ab[0][6] ));
   NOR2 \mult_20_3/AN1_0_5  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [5]),
	.OUT(\mult_20_3/ab[0][5] ));
   NOR2 \mult_20_3/AN1_0_4  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [4]),
	.OUT(\mult_20_3/ab[0][4] ));
   NOR2 \mult_20_3/AN1_0_3  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [3]),
	.OUT(\mult_20_3/ab[0][3] ));
   NOR2 \mult_20_3/AN1_0_2  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [2]),
	.OUT(\mult_20_3/ab[0][2] ));
   NOR2 \mult_20_3/AN1_0_1  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [1]),
	.OUT(\mult_20_3/ab[0][1] ));
   NOR2 \mult_20_3/AN1_0_0_0  (.A(\mult_20_3/A_notx [0]),
	.B(\mult_20_3/B_notx [0]),
	.OUT(N129));
   OAI21 \mult_20_2/FS_1/U6_1_0_3  (.OUT(\mult_20_2/FS_1/C[1][3][0] ),
	.C(n3129),
	.B(n3128),
	.A(n3127));
   OAI21 \mult_20_2/FS_1/U6_0_3_1  (.OUT(\mult_20_2/FS_1/C[1][3][1] ),
	.C(\mult_20_2/FS_1/G_n_int[0][3][0] ),
	.B(n3125),
	.A(n3124));
   XOR2 \mult_20_2/FS_1/U3_C_0_3_1  (.A(\mult_20_2/FS_1/PG_int[0][3][1] ),
	.B(\mult_20_2/FS_1/C[1][3][1] ),
	.OUT(N112));
   XOR2 \mult_20_2/FS_1/U3_C_0_3_0  (.A(\mult_20_2/FS_1/PG_int[0][3][0] ),
	.B(\mult_20_2/FS_1/C[1][3][0] ),
	.OUT(N111));
   NAND2 \mult_20_2/FS_1/U3_B_0_3_0  (.A(\mult_20_2/FS_1/G_n_int[0][3][0] ),
	.B(\mult_20_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3121));
   NAND2 \mult_20_2/FS_1/U2_0_3_0  (.A(\mult_20_2/A1[12] ),
	.B(\mult_20_2/A2[12] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_20_2/FS_1/U1_0_3_0  (.A(n3119),
	.B(n3120),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_20_2/FS_1/U6_0_2_3  (.OUT(\mult_20_2/FS_1/C[1][2][3] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][2] ),
	.B(n3118),
	.A(n3117));
   OAI21 \mult_20_2/FS_1/U5_0_2_3  (.OUT(\mult_20_2/FS_1/G[1][0][2] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][3] ),
	.B(n3116),
	.A(n3115));
   NAND2 \mult_20_2/FS_1/U4_0_2_3  (.A(\mult_20_2/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_20_2/FS_1/P[0][2][3] ),
	.OUT(n3128));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_3  (.A(\mult_20_2/FS_1/PG_int[0][2][3] ),
	.B(\mult_20_2/FS_1/C[1][2][3] ),
	.OUT(N110));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_3  (.A(\mult_20_2/FS_1/G_n_int[0][2][3] ),
	.B(\mult_20_2/FS_1/P[0][2][3] ),
	.OUT(n3114));
   NAND2 \mult_20_2/FS_1/U2_0_2_3  (.A(\mult_20_2/A1[11] ),
	.B(\mult_20_2/A2[11] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_3  (.A(n3112),
	.B(n3113),
	.OUT(\mult_20_2/FS_1/P[0][2][3] ));
   OAI21 \mult_20_2/FS_1/U6_0_2_2  (.OUT(\mult_20_2/FS_1/C[1][2][2] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][1] ),
	.B(n3111),
	.A(n3110));
   OAI21 \mult_20_2/FS_1/U5_0_2_2  (.OUT(\mult_20_2/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][2] ),
	.B(n3118),
	.A(n3109));
   NAND2 \mult_20_2/FS_1/U4_0_2_2  (.A(\mult_20_2/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_20_2/FS_1/P[0][2][2] ),
	.OUT(n3108));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_2  (.A(\mult_20_2/FS_1/PG_int[0][2][2] ),
	.B(\mult_20_2/FS_1/C[1][2][2] ),
	.OUT(N109));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_2  (.A(\mult_20_2/FS_1/G_n_int[0][2][2] ),
	.B(\mult_20_2/FS_1/P[0][2][2] ),
	.OUT(n3107));
   NAND2 \mult_20_2/FS_1/U2_0_2_2  (.A(\mult_20_2/A1[10] ),
	.B(\mult_20_2/A2[10] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_2  (.A(n3105),
	.B(n3106),
	.OUT(\mult_20_2/FS_1/P[0][2][2] ));
   OAI21 \mult_20_2/FS_1/U6_0_2_1  (.OUT(\mult_20_2/FS_1/C[1][2][1] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][0] ),
	.B(n3104),
	.A(n3127));
   OAI21 \mult_20_2/FS_1/U5_0_2_1  (.OUT(\mult_20_2/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_20_2/FS_1/G_n_int[0][2][1] ),
	.B(n3111),
	.A(\mult_20_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_2/FS_1/U4_0_2_1  (.A(\mult_20_2/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_20_2/FS_1/P[0][2][1] ),
	.OUT(n3103));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_1  (.A(\mult_20_2/FS_1/PG_int[0][2][1] ),
	.B(\mult_20_2/FS_1/C[1][2][1] ),
	.OUT(N108));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_1  (.A(\mult_20_2/FS_1/G_n_int[0][2][1] ),
	.B(\mult_20_2/FS_1/P[0][2][1] ),
	.OUT(n3102));
   NAND2 \mult_20_2/FS_1/U2_0_2_1  (.A(\mult_20_2/A1[9] ),
	.B(\mult_20_2/A2[9] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_1  (.A(n3100),
	.B(n3101),
	.OUT(\mult_20_2/FS_1/P[0][2][1] ));
   XOR2 \mult_20_2/FS_1/U3_C_0_2_0  (.A(\mult_20_2/FS_1/PG_int[0][2][0] ),
	.B(\mult_20_2/FS_1/C[1][2][0] ),
	.OUT(N107));
   NAND2 \mult_20_2/FS_1/U3_B_0_2_0  (.A(\mult_20_2/FS_1/G_n_int[0][2][0] ),
	.B(\mult_20_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3099));
   NAND2 \mult_20_2/FS_1/U2_0_2_0  (.A(\mult_20_2/A1[8] ),
	.B(\mult_20_2/A2[8] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20_2/FS_1/U1_0_2_0  (.A(n3097),
	.B(n3098),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_20_2/FS_1/U3_B_0_1_3  (.A(\mult_20_2/FS_1/G_n_int[0][1][3] ),
	.B(\mult_20_2/FS_1/P[0][1][3] ),
	.OUT(n3096));
   NAND2 \mult_20_2/FS_1/U2_0_1_3  (.A(\mult_20_2/A1[7] ),
	.B(\mult_20_2/A2[7] ),
	.OUT(\mult_20_2/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_20_2/FS_1/U1_0_1_3  (.A(n3094),
	.B(n3095),
	.OUT(\mult_20_2/FS_1/P[0][1][3] ));
   INVERTER \mult_20_2/AN1_7  (.IN(matrix11[7]),
	.OUT(\mult_20_2/A_not[7] ));
   INVERTER \mult_20_2/AN1_6  (.IN(matrix11[6]),
	.OUT(\mult_20_2/A_notx [6]));
   INVERTER \mult_20_2/AN1_5  (.IN(matrix11[5]),
	.OUT(\mult_20_2/A_notx [5]));
   INVERTER \mult_20_2/AN1_4  (.IN(matrix11[4]),
	.OUT(\mult_20_2/A_notx [4]));
   INVERTER \mult_20_2/AN1_3  (.IN(matrix11[3]),
	.OUT(\mult_20_2/A_notx [3]));
   INVERTER \mult_20_2/AN1_2  (.IN(matrix11[2]),
	.OUT(\mult_20_2/A_notx [2]));
   INVERTER \mult_20_2/AN1_1  (.IN(matrix11[1]),
	.OUT(\mult_20_2/A_notx [1]));
   INVERTER \mult_20_2/AN1_0  (.IN(matrix11[0]),
	.OUT(\mult_20_2/A_notx [0]));
   INVERTER \mult_20_2/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_20_2/B_not[7] ));
   INVERTER \mult_20_2/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_20_2/B_notx [6]));
   INVERTER \mult_20_2/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_20_2/B_notx [5]));
   INVERTER \mult_20_2/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_20_2/B_notx [4]));
   INVERTER \mult_20_2/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_20_2/B_notx [3]));
   INVERTER \mult_20_2/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_20_2/B_notx [2]));
   INVERTER \mult_20_2/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_20_2/B_notx [1]));
   INVERTER \mult_20_2/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_20_2/B_notx [0]));
   NOR2 \mult_20_2/AN1_7_7  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[7][7] ));
   NOR2 \mult_20_2/AN3_7_6  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[7][6] ));
   NOR2 \mult_20_2/AN3_7_5  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[7][5] ));
   NOR2 \mult_20_2/AN3_7_4  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[7][4] ));
   NOR2 \mult_20_2/AN3_7_3  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[7][3] ));
   NOR2 \mult_20_2/AN3_7_2  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[7][2] ));
   NOR2 \mult_20_2/AN3_7_1  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[7][1] ));
   NOR2 \mult_20_2/AN3_7_0  (.A(\mult_20_2/A_not[7] ),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[7][0] ));
   NOR2 \mult_20_2/AN2_6_7  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[6][7] ));
   NOR2 \mult_20_2/AN1_6_6  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[6][6] ));
   NOR2 \mult_20_2/AN1_6_5  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[6][5] ));
   NOR2 \mult_20_2/AN1_6_4  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[6][4] ));
   NOR2 \mult_20_2/AN1_6_3  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[6][3] ));
   NOR2 \mult_20_2/AN1_6_2  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[6][2] ));
   NOR2 \mult_20_2/AN1_6_1  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[6][1] ));
   NOR2 \mult_20_2/AN1_6_0_0  (.A(\mult_20_2/A_notx [6]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[6][0] ));
   NOR2 \mult_20_2/AN2_5_7  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[5][7] ));
   NOR2 \mult_20_2/AN1_5_6  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[5][6] ));
   NOR2 \mult_20_2/AN1_5_5  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[5][5] ));
   NOR2 \mult_20_2/AN1_5_4  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[5][4] ));
   NOR2 \mult_20_2/AN1_5_3  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[5][3] ));
   NOR2 \mult_20_2/AN1_5_2  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[5][2] ));
   NOR2 \mult_20_2/AN1_5_1  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[5][1] ));
   NOR2 \mult_20_2/AN1_5_0_0  (.A(\mult_20_2/A_notx [5]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[5][0] ));
   NOR2 \mult_20_2/AN2_4_7  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[4][7] ));
   NOR2 \mult_20_2/AN1_4_6  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[4][6] ));
   NOR2 \mult_20_2/AN1_4_5  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[4][5] ));
   NOR2 \mult_20_2/AN1_4_4  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[4][4] ));
   NOR2 \mult_20_2/AN1_4_3  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[4][3] ));
   NOR2 \mult_20_2/AN1_4_2  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[4][2] ));
   NOR2 \mult_20_2/AN1_4_1  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[4][1] ));
   NOR2 \mult_20_2/AN1_4_0_0  (.A(\mult_20_2/A_notx [4]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[4][0] ));
   NOR2 \mult_20_2/AN2_3_7  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[3][7] ));
   NOR2 \mult_20_2/AN1_3_6  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[3][6] ));
   NOR2 \mult_20_2/AN1_3_5  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[3][5] ));
   NOR2 \mult_20_2/AN1_3_4  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[3][4] ));
   NOR2 \mult_20_2/AN1_3_3  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[3][3] ));
   NOR2 \mult_20_2/AN1_3_2  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[3][2] ));
   NOR2 \mult_20_2/AN1_3_1  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[3][1] ));
   NOR2 \mult_20_2/AN1_3_0_0  (.A(\mult_20_2/A_notx [3]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[3][0] ));
   NOR2 \mult_20_2/AN2_2_7  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[2][7] ));
   NOR2 \mult_20_2/AN1_2_6  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[2][6] ));
   NOR2 \mult_20_2/AN1_2_5  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[2][5] ));
   NOR2 \mult_20_2/AN1_2_4  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[2][4] ));
   NOR2 \mult_20_2/AN1_2_3  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[2][3] ));
   NOR2 \mult_20_2/AN1_2_2  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[2][2] ));
   NOR2 \mult_20_2/AN1_2_1  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[2][1] ));
   NOR2 \mult_20_2/AN1_2_0_0  (.A(\mult_20_2/A_notx [2]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[2][0] ));
   NOR2 \mult_20_2/AN2_1_7  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[1][7] ));
   NOR2 \mult_20_2/AN1_1_6  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[1][6] ));
   NOR2 \mult_20_2/AN1_1_5  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[1][5] ));
   NOR2 \mult_20_2/AN1_1_4  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[1][4] ));
   NOR2 \mult_20_2/AN1_1_3  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[1][3] ));
   NOR2 \mult_20_2/AN1_1_2  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[1][2] ));
   NOR2 \mult_20_2/AN1_1_1  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[1][1] ));
   NOR2 \mult_20_2/AN1_1_0_0  (.A(\mult_20_2/A_notx [1]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(\mult_20_2/ab[1][0] ));
   NOR2 \mult_20_2/AN2_0_7  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_not[7] ),
	.OUT(\mult_20_2/ab[0][7] ));
   NOR2 \mult_20_2/AN1_0_6  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [6]),
	.OUT(\mult_20_2/ab[0][6] ));
   NOR2 \mult_20_2/AN1_0_5  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [5]),
	.OUT(\mult_20_2/ab[0][5] ));
   NOR2 \mult_20_2/AN1_0_4  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [4]),
	.OUT(\mult_20_2/ab[0][4] ));
   NOR2 \mult_20_2/AN1_0_3  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [3]),
	.OUT(\mult_20_2/ab[0][3] ));
   NOR2 \mult_20_2/AN1_0_2  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [2]),
	.OUT(\mult_20_2/ab[0][2] ));
   NOR2 \mult_20_2/AN1_0_1  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [1]),
	.OUT(\mult_20_2/ab[0][1] ));
   NOR2 \mult_20_2/AN1_0_0_0  (.A(\mult_20_2/A_notx [0]),
	.B(\mult_20_2/B_notx [0]),
	.OUT(N97));
   OAI21 \mult_20/FS_1/U6_1_0_3  (.OUT(\mult_20/FS_1/C[1][3][0] ),
	.C(n3079),
	.B(n3078),
	.A(n3077));
   OAI21 \mult_20/FS_1/U6_0_3_1  (.OUT(\mult_20/FS_1/C[1][3][1] ),
	.C(\mult_20/FS_1/G_n_int[0][3][0] ),
	.B(n3075),
	.A(n3074));
   XOR2 \mult_20/FS_1/U3_C_0_3_1  (.A(\mult_20/FS_1/PG_int[0][3][1] ),
	.B(\mult_20/FS_1/C[1][3][1] ),
	.OUT(N96));
   XOR2 \mult_20/FS_1/U3_C_0_3_0  (.A(\mult_20/FS_1/PG_int[0][3][0] ),
	.B(\mult_20/FS_1/C[1][3][0] ),
	.OUT(N95));
   NAND2 \mult_20/FS_1/U3_B_0_3_0  (.A(\mult_20/FS_1/G_n_int[0][3][0] ),
	.B(\mult_20/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3071));
   NAND2 \mult_20/FS_1/U2_0_3_0  (.A(\mult_20/A1[12] ),
	.B(\mult_20/A2[12] ),
	.OUT(\mult_20/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_20/FS_1/U1_0_3_0  (.A(n3069),
	.B(n3070),
	.OUT(\mult_20/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_20/FS_1/U6_0_2_3  (.OUT(\mult_20/FS_1/C[1][2][3] ),
	.C(\mult_20/FS_1/G_n_int[0][2][2] ),
	.B(n3068),
	.A(n3067));
   OAI21 \mult_20/FS_1/U5_0_2_3  (.OUT(\mult_20/FS_1/G[1][0][2] ),
	.C(\mult_20/FS_1/G_n_int[0][2][3] ),
	.B(n3066),
	.A(n3065));
   NAND2 \mult_20/FS_1/U4_0_2_3  (.A(\mult_20/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_20/FS_1/P[0][2][3] ),
	.OUT(n3078));
   XOR2 \mult_20/FS_1/U3_C_0_2_3  (.A(\mult_20/FS_1/PG_int[0][2][3] ),
	.B(\mult_20/FS_1/C[1][2][3] ),
	.OUT(N94));
   NAND2 \mult_20/FS_1/U3_B_0_2_3  (.A(\mult_20/FS_1/G_n_int[0][2][3] ),
	.B(\mult_20/FS_1/P[0][2][3] ),
	.OUT(n3064));
   NAND2 \mult_20/FS_1/U2_0_2_3  (.A(\mult_20/A1[11] ),
	.B(\mult_20/A2[11] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_20/FS_1/U1_0_2_3  (.A(n3062),
	.B(n3063),
	.OUT(\mult_20/FS_1/P[0][2][3] ));
   OAI21 \mult_20/FS_1/U6_0_2_2  (.OUT(\mult_20/FS_1/C[1][2][2] ),
	.C(\mult_20/FS_1/G_n_int[0][2][1] ),
	.B(n3061),
	.A(n3060));
   OAI21 \mult_20/FS_1/U5_0_2_2  (.OUT(\mult_20/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_20/FS_1/G_n_int[0][2][2] ),
	.B(n3068),
	.A(n3059));
   NAND2 \mult_20/FS_1/U4_0_2_2  (.A(\mult_20/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_20/FS_1/P[0][2][2] ),
	.OUT(n3058));
   XOR2 \mult_20/FS_1/U3_C_0_2_2  (.A(\mult_20/FS_1/PG_int[0][2][2] ),
	.B(\mult_20/FS_1/C[1][2][2] ),
	.OUT(N93));
   NAND2 \mult_20/FS_1/U3_B_0_2_2  (.A(\mult_20/FS_1/G_n_int[0][2][2] ),
	.B(\mult_20/FS_1/P[0][2][2] ),
	.OUT(n3057));
   NAND2 \mult_20/FS_1/U2_0_2_2  (.A(\mult_20/A1[10] ),
	.B(\mult_20/A2[10] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_20/FS_1/U1_0_2_2  (.A(n3055),
	.B(n3056),
	.OUT(\mult_20/FS_1/P[0][2][2] ));
   OAI21 \mult_20/FS_1/U6_0_2_1  (.OUT(\mult_20/FS_1/C[1][2][1] ),
	.C(\mult_20/FS_1/G_n_int[0][2][0] ),
	.B(n3054),
	.A(n3077));
   OAI21 \mult_20/FS_1/U5_0_2_1  (.OUT(\mult_20/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_20/FS_1/G_n_int[0][2][1] ),
	.B(n3061),
	.A(\mult_20/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20/FS_1/U4_0_2_1  (.A(\mult_20/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_20/FS_1/P[0][2][1] ),
	.OUT(n3053));
   XOR2 \mult_20/FS_1/U3_C_0_2_1  (.A(\mult_20/FS_1/PG_int[0][2][1] ),
	.B(\mult_20/FS_1/C[1][2][1] ),
	.OUT(N92));
   NAND2 \mult_20/FS_1/U3_B_0_2_1  (.A(\mult_20/FS_1/G_n_int[0][2][1] ),
	.B(\mult_20/FS_1/P[0][2][1] ),
	.OUT(n3052));
   NAND2 \mult_20/FS_1/U2_0_2_1  (.A(\mult_20/A1[9] ),
	.B(\mult_20/A2[9] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_20/FS_1/U1_0_2_1  (.A(n3050),
	.B(n3051),
	.OUT(\mult_20/FS_1/P[0][2][1] ));
   XOR2 \mult_20/FS_1/U3_C_0_2_0  (.A(\mult_20/FS_1/PG_int[0][2][0] ),
	.B(\mult_20/FS_1/C[1][2][0] ),
	.OUT(N91));
   NAND2 \mult_20/FS_1/U3_B_0_2_0  (.A(\mult_20/FS_1/G_n_int[0][2][0] ),
	.B(\mult_20/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3049));
   NAND2 \mult_20/FS_1/U2_0_2_0  (.A(\mult_20/A1[8] ),
	.B(\mult_20/A2[8] ),
	.OUT(\mult_20/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_20/FS_1/U1_0_2_0  (.A(n3047),
	.B(n3048),
	.OUT(\mult_20/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_20/FS_1/U3_B_0_1_3  (.A(\mult_20/FS_1/G_n_int[0][1][3] ),
	.B(\mult_20/FS_1/P[0][1][3] ),
	.OUT(n3046));
   NAND2 \mult_20/FS_1/U2_0_1_3  (.A(\mult_20/A1[7] ),
	.B(\mult_20/A2[7] ),
	.OUT(\mult_20/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_20/FS_1/U1_0_1_3  (.A(n3044),
	.B(n3045),
	.OUT(\mult_20/FS_1/P[0][1][3] ));
   INVERTER \mult_20/AN1_7  (.IN(matrix10[7]),
	.OUT(\mult_20/A_not[7] ));
   INVERTER \mult_20/AN1_6  (.IN(matrix10[6]),
	.OUT(\mult_20/A_notx [6]));
   INVERTER \mult_20/AN1_5  (.IN(matrix10[5]),
	.OUT(\mult_20/A_notx [5]));
   INVERTER \mult_20/AN1_4  (.IN(matrix10[4]),
	.OUT(\mult_20/A_notx [4]));
   INVERTER \mult_20/AN1_3  (.IN(matrix10[3]),
	.OUT(\mult_20/A_notx [3]));
   INVERTER \mult_20/AN1_2  (.IN(matrix10[2]),
	.OUT(\mult_20/A_notx [2]));
   INVERTER \mult_20/AN1_1  (.IN(matrix10[1]),
	.OUT(\mult_20/A_notx [1]));
   INVERTER \mult_20/AN1_0  (.IN(matrix10[0]),
	.OUT(\mult_20/A_notx [0]));
   INVERTER \mult_20/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_20/B_not[7] ));
   INVERTER \mult_20/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_20/B_notx [6]));
   INVERTER \mult_20/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_20/B_notx [5]));
   INVERTER \mult_20/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_20/B_notx [4]));
   INVERTER \mult_20/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_20/B_notx [3]));
   INVERTER \mult_20/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_20/B_notx [2]));
   INVERTER \mult_20/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_20/B_notx [1]));
   INVERTER \mult_20/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_20/B_notx [0]));
   NOR2 \mult_20/AN1_7_7  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[7][7] ));
   NOR2 \mult_20/AN3_7_6  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[7][6] ));
   NOR2 \mult_20/AN3_7_5  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[7][5] ));
   NOR2 \mult_20/AN3_7_4  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[7][4] ));
   NOR2 \mult_20/AN3_7_3  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[7][3] ));
   NOR2 \mult_20/AN3_7_2  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[7][2] ));
   NOR2 \mult_20/AN3_7_1  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[7][1] ));
   NOR2 \mult_20/AN3_7_0  (.A(\mult_20/A_not[7] ),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[7][0] ));
   NOR2 \mult_20/AN2_6_7  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[6][7] ));
   NOR2 \mult_20/AN1_6_6  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[6][6] ));
   NOR2 \mult_20/AN1_6_5  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[6][5] ));
   NOR2 \mult_20/AN1_6_4  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[6][4] ));
   NOR2 \mult_20/AN1_6_3  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[6][3] ));
   NOR2 \mult_20/AN1_6_2  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[6][2] ));
   NOR2 \mult_20/AN1_6_1  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[6][1] ));
   NOR2 \mult_20/AN1_6_0_0  (.A(\mult_20/A_notx [6]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[6][0] ));
   NOR2 \mult_20/AN2_5_7  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[5][7] ));
   NOR2 \mult_20/AN1_5_6  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[5][6] ));
   NOR2 \mult_20/AN1_5_5  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[5][5] ));
   NOR2 \mult_20/AN1_5_4  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[5][4] ));
   NOR2 \mult_20/AN1_5_3  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[5][3] ));
   NOR2 \mult_20/AN1_5_2  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[5][2] ));
   NOR2 \mult_20/AN1_5_1  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[5][1] ));
   NOR2 \mult_20/AN1_5_0_0  (.A(\mult_20/A_notx [5]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[5][0] ));
   NOR2 \mult_20/AN2_4_7  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[4][7] ));
   NOR2 \mult_20/AN1_4_6  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[4][6] ));
   NOR2 \mult_20/AN1_4_5  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[4][5] ));
   NOR2 \mult_20/AN1_4_4  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[4][4] ));
   NOR2 \mult_20/AN1_4_3  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[4][3] ));
   NOR2 \mult_20/AN1_4_2  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[4][2] ));
   NOR2 \mult_20/AN1_4_1  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[4][1] ));
   NOR2 \mult_20/AN1_4_0_0  (.A(\mult_20/A_notx [4]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[4][0] ));
   NOR2 \mult_20/AN2_3_7  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[3][7] ));
   NOR2 \mult_20/AN1_3_6  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[3][6] ));
   NOR2 \mult_20/AN1_3_5  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[3][5] ));
   NOR2 \mult_20/AN1_3_4  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[3][4] ));
   NOR2 \mult_20/AN1_3_3  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[3][3] ));
   NOR2 \mult_20/AN1_3_2  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[3][2] ));
   NOR2 \mult_20/AN1_3_1  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[3][1] ));
   NOR2 \mult_20/AN1_3_0_0  (.A(\mult_20/A_notx [3]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[3][0] ));
   NOR2 \mult_20/AN2_2_7  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[2][7] ));
   NOR2 \mult_20/AN1_2_6  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[2][6] ));
   NOR2 \mult_20/AN1_2_5  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[2][5] ));
   NOR2 \mult_20/AN1_2_4  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[2][4] ));
   NOR2 \mult_20/AN1_2_3  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[2][3] ));
   NOR2 \mult_20/AN1_2_2  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[2][2] ));
   NOR2 \mult_20/AN1_2_1  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[2][1] ));
   NOR2 \mult_20/AN1_2_0_0  (.A(\mult_20/A_notx [2]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[2][0] ));
   NOR2 \mult_20/AN2_1_7  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[1][7] ));
   NOR2 \mult_20/AN1_1_6  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[1][6] ));
   NOR2 \mult_20/AN1_1_5  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[1][5] ));
   NOR2 \mult_20/AN1_1_4  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[1][4] ));
   NOR2 \mult_20/AN1_1_3  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[1][3] ));
   NOR2 \mult_20/AN1_1_2  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[1][2] ));
   NOR2 \mult_20/AN1_1_1  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[1][1] ));
   NOR2 \mult_20/AN1_1_0_0  (.A(\mult_20/A_notx [1]),
	.B(\mult_20/B_notx [0]),
	.OUT(\mult_20/ab[1][0] ));
   NOR2 \mult_20/AN2_0_7  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_not[7] ),
	.OUT(\mult_20/ab[0][7] ));
   NOR2 \mult_20/AN1_0_6  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [6]),
	.OUT(\mult_20/ab[0][6] ));
   NOR2 \mult_20/AN1_0_5  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [5]),
	.OUT(\mult_20/ab[0][5] ));
   NOR2 \mult_20/AN1_0_4  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [4]),
	.OUT(\mult_20/ab[0][4] ));
   NOR2 \mult_20/AN1_0_3  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [3]),
	.OUT(\mult_20/ab[0][3] ));
   NOR2 \mult_20/AN1_0_2  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [2]),
	.OUT(\mult_20/ab[0][2] ));
   NOR2 \mult_20/AN1_0_1  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [1]),
	.OUT(\mult_20/ab[0][1] ));
   NOR2 \mult_20/AN1_0_0_0  (.A(\mult_20/A_notx [0]),
	.B(\mult_20/B_notx [0]),
	.OUT(N81));
   OAI21 \mult_19_3/FS_1/U6_1_0_3  (.OUT(\mult_19_3/FS_1/C[1][3][0] ),
	.C(n3029),
	.B(n3028),
	.A(n3027));
   OAI21 \mult_19_3/FS_1/U6_0_3_1  (.OUT(\mult_19_3/FS_1/C[1][3][1] ),
	.C(\mult_19_3/FS_1/G_n_int[0][3][0] ),
	.B(n3025),
	.A(n3024));
   XOR2 \mult_19_3/FS_1/U3_C_0_3_1  (.A(\mult_19_3/FS_1/PG_int[0][3][1] ),
	.B(\mult_19_3/FS_1/C[1][3][1] ),
	.OUT(N64));
   XOR2 \mult_19_3/FS_1/U3_C_0_3_0  (.A(\mult_19_3/FS_1/PG_int[0][3][0] ),
	.B(\mult_19_3/FS_1/C[1][3][0] ),
	.OUT(N63));
   NAND2 \mult_19_3/FS_1/U3_B_0_3_0  (.A(\mult_19_3/FS_1/G_n_int[0][3][0] ),
	.B(\mult_19_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3021));
   NAND2 \mult_19_3/FS_1/U2_0_3_0  (.A(\mult_19_3/A1[12] ),
	.B(\mult_19_3/A2[12] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_19_3/FS_1/U1_0_3_0  (.A(n3019),
	.B(n3020),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_19_3/FS_1/U6_0_2_3  (.OUT(\mult_19_3/FS_1/C[1][2][3] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][2] ),
	.B(n3018),
	.A(n3017));
   OAI21 \mult_19_3/FS_1/U5_0_2_3  (.OUT(\mult_19_3/FS_1/G[1][0][2] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][3] ),
	.B(n3016),
	.A(n3015));
   NAND2 \mult_19_3/FS_1/U4_0_2_3  (.A(\mult_19_3/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_19_3/FS_1/P[0][2][3] ),
	.OUT(n3028));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_3  (.A(\mult_19_3/FS_1/PG_int[0][2][3] ),
	.B(\mult_19_3/FS_1/C[1][2][3] ),
	.OUT(N62));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_3  (.A(\mult_19_3/FS_1/G_n_int[0][2][3] ),
	.B(\mult_19_3/FS_1/P[0][2][3] ),
	.OUT(n3014));
   NAND2 \mult_19_3/FS_1/U2_0_2_3  (.A(\mult_19_3/A1[11] ),
	.B(\mult_19_3/A2[11] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_3  (.A(n3012),
	.B(n3013),
	.OUT(\mult_19_3/FS_1/P[0][2][3] ));
   OAI21 \mult_19_3/FS_1/U6_0_2_2  (.OUT(\mult_19_3/FS_1/C[1][2][2] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][1] ),
	.B(n3011),
	.A(n3010));
   OAI21 \mult_19_3/FS_1/U5_0_2_2  (.OUT(\mult_19_3/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][2] ),
	.B(n3018),
	.A(n3009));
   NAND2 \mult_19_3/FS_1/U4_0_2_2  (.A(\mult_19_3/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_19_3/FS_1/P[0][2][2] ),
	.OUT(n3008));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_2  (.A(\mult_19_3/FS_1/PG_int[0][2][2] ),
	.B(\mult_19_3/FS_1/C[1][2][2] ),
	.OUT(N61));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_2  (.A(\mult_19_3/FS_1/G_n_int[0][2][2] ),
	.B(\mult_19_3/FS_1/P[0][2][2] ),
	.OUT(n3007));
   NAND2 \mult_19_3/FS_1/U2_0_2_2  (.A(\mult_19_3/A1[10] ),
	.B(\mult_19_3/A2[10] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_2  (.A(n3005),
	.B(n3006),
	.OUT(\mult_19_3/FS_1/P[0][2][2] ));
   OAI21 \mult_19_3/FS_1/U6_0_2_1  (.OUT(\mult_19_3/FS_1/C[1][2][1] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][0] ),
	.B(n3004),
	.A(n3027));
   OAI21 \mult_19_3/FS_1/U5_0_2_1  (.OUT(\mult_19_3/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_19_3/FS_1/G_n_int[0][2][1] ),
	.B(n3011),
	.A(\mult_19_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_3/FS_1/U4_0_2_1  (.A(\mult_19_3/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_19_3/FS_1/P[0][2][1] ),
	.OUT(n3003));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_1  (.A(\mult_19_3/FS_1/PG_int[0][2][1] ),
	.B(\mult_19_3/FS_1/C[1][2][1] ),
	.OUT(N60));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_1  (.A(\mult_19_3/FS_1/G_n_int[0][2][1] ),
	.B(\mult_19_3/FS_1/P[0][2][1] ),
	.OUT(n3002));
   NAND2 \mult_19_3/FS_1/U2_0_2_1  (.A(\mult_19_3/A1[9] ),
	.B(\mult_19_3/A2[9] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_1  (.A(n3000),
	.B(n3001),
	.OUT(\mult_19_3/FS_1/P[0][2][1] ));
   XOR2 \mult_19_3/FS_1/U3_C_0_2_0  (.A(\mult_19_3/FS_1/PG_int[0][2][0] ),
	.B(\mult_19_3/FS_1/C[1][2][0] ),
	.OUT(N59));
   NAND2 \mult_19_3/FS_1/U3_B_0_2_0  (.A(\mult_19_3/FS_1/G_n_int[0][2][0] ),
	.B(\mult_19_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2999));
   NAND2 \mult_19_3/FS_1/U2_0_2_0  (.A(\mult_19_3/A1[8] ),
	.B(\mult_19_3/A2[8] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_3/FS_1/U1_0_2_0  (.A(n2997),
	.B(n2998),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_19_3/FS_1/U3_B_0_1_3  (.A(\mult_19_3/FS_1/G_n_int[0][1][3] ),
	.B(\mult_19_3/FS_1/P[0][1][3] ),
	.OUT(n2996));
   NAND2 \mult_19_3/FS_1/U2_0_1_3  (.A(\mult_19_3/A1[7] ),
	.B(\mult_19_3/A2[7] ),
	.OUT(\mult_19_3/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_19_3/FS_1/U1_0_1_3  (.A(n2994),
	.B(n2995),
	.OUT(\mult_19_3/FS_1/P[0][1][3] ));
   INVERTER \mult_19_3/AN1_7  (.IN(matrix02[7]),
	.OUT(\mult_19_3/A_not[7] ));
   INVERTER \mult_19_3/AN1_6  (.IN(matrix02[6]),
	.OUT(\mult_19_3/A_notx [6]));
   INVERTER \mult_19_3/AN1_5  (.IN(matrix02[5]),
	.OUT(\mult_19_3/A_notx [5]));
   INVERTER \mult_19_3/AN1_4  (.IN(matrix02[4]),
	.OUT(\mult_19_3/A_notx [4]));
   INVERTER \mult_19_3/AN1_3  (.IN(matrix02[3]),
	.OUT(\mult_19_3/A_notx [3]));
   INVERTER \mult_19_3/AN1_2  (.IN(matrix02[2]),
	.OUT(\mult_19_3/A_notx [2]));
   INVERTER \mult_19_3/AN1_1  (.IN(matrix02[1]),
	.OUT(\mult_19_3/A_notx [1]));
   INVERTER \mult_19_3/AN1_0  (.IN(matrix02[0]),
	.OUT(\mult_19_3/A_notx [0]));
   INVERTER \mult_19_3/AN1_7_0  (.IN(vector_2[7]),
	.OUT(\mult_19_3/B_not[7] ));
   INVERTER \mult_19_3/AN1_6_0  (.IN(vector_2[6]),
	.OUT(\mult_19_3/B_notx [6]));
   INVERTER \mult_19_3/AN1_5_0  (.IN(vector_2[5]),
	.OUT(\mult_19_3/B_notx [5]));
   INVERTER \mult_19_3/AN1_4_0  (.IN(vector_2[4]),
	.OUT(\mult_19_3/B_notx [4]));
   INVERTER \mult_19_3/AN1_3_0  (.IN(vector_2[3]),
	.OUT(\mult_19_3/B_notx [3]));
   INVERTER \mult_19_3/AN1_2_0  (.IN(vector_2[2]),
	.OUT(\mult_19_3/B_notx [2]));
   INVERTER \mult_19_3/AN1_1_0  (.IN(vector_2[1]),
	.OUT(\mult_19_3/B_notx [1]));
   INVERTER \mult_19_3/AN1_0_0  (.IN(vector_2[0]),
	.OUT(\mult_19_3/B_notx [0]));
   NOR2 \mult_19_3/AN1_7_7  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[7][7] ));
   NOR2 \mult_19_3/AN3_7_6  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[7][6] ));
   NOR2 \mult_19_3/AN3_7_5  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[7][5] ));
   NOR2 \mult_19_3/AN3_7_4  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[7][4] ));
   NOR2 \mult_19_3/AN3_7_3  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[7][3] ));
   NOR2 \mult_19_3/AN3_7_2  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[7][2] ));
   NOR2 \mult_19_3/AN3_7_1  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[7][1] ));
   NOR2 \mult_19_3/AN3_7_0  (.A(\mult_19_3/A_not[7] ),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[7][0] ));
   NOR2 \mult_19_3/AN2_6_7  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[6][7] ));
   NOR2 \mult_19_3/AN1_6_6  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[6][6] ));
   NOR2 \mult_19_3/AN1_6_5  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[6][5] ));
   NOR2 \mult_19_3/AN1_6_4  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[6][4] ));
   NOR2 \mult_19_3/AN1_6_3  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[6][3] ));
   NOR2 \mult_19_3/AN1_6_2  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[6][2] ));
   NOR2 \mult_19_3/AN1_6_1  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[6][1] ));
   NOR2 \mult_19_3/AN1_6_0_0  (.A(\mult_19_3/A_notx [6]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[6][0] ));
   NOR2 \mult_19_3/AN2_5_7  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[5][7] ));
   NOR2 \mult_19_3/AN1_5_6  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[5][6] ));
   NOR2 \mult_19_3/AN1_5_5  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[5][5] ));
   NOR2 \mult_19_3/AN1_5_4  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[5][4] ));
   NOR2 \mult_19_3/AN1_5_3  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[5][3] ));
   NOR2 \mult_19_3/AN1_5_2  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[5][2] ));
   NOR2 \mult_19_3/AN1_5_1  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[5][1] ));
   NOR2 \mult_19_3/AN1_5_0_0  (.A(\mult_19_3/A_notx [5]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[5][0] ));
   NOR2 \mult_19_3/AN2_4_7  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[4][7] ));
   NOR2 \mult_19_3/AN1_4_6  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[4][6] ));
   NOR2 \mult_19_3/AN1_4_5  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[4][5] ));
   NOR2 \mult_19_3/AN1_4_4  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[4][4] ));
   NOR2 \mult_19_3/AN1_4_3  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[4][3] ));
   NOR2 \mult_19_3/AN1_4_2  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[4][2] ));
   NOR2 \mult_19_3/AN1_4_1  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[4][1] ));
   NOR2 \mult_19_3/AN1_4_0_0  (.A(\mult_19_3/A_notx [4]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[4][0] ));
   NOR2 \mult_19_3/AN2_3_7  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[3][7] ));
   NOR2 \mult_19_3/AN1_3_6  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[3][6] ));
   NOR2 \mult_19_3/AN1_3_5  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[3][5] ));
   NOR2 \mult_19_3/AN1_3_4  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[3][4] ));
   NOR2 \mult_19_3/AN1_3_3  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[3][3] ));
   NOR2 \mult_19_3/AN1_3_2  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[3][2] ));
   NOR2 \mult_19_3/AN1_3_1  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[3][1] ));
   NOR2 \mult_19_3/AN1_3_0_0  (.A(\mult_19_3/A_notx [3]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[3][0] ));
   NOR2 \mult_19_3/AN2_2_7  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[2][7] ));
   NOR2 \mult_19_3/AN1_2_6  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[2][6] ));
   NOR2 \mult_19_3/AN1_2_5  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[2][5] ));
   NOR2 \mult_19_3/AN1_2_4  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[2][4] ));
   NOR2 \mult_19_3/AN1_2_3  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[2][3] ));
   NOR2 \mult_19_3/AN1_2_2  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[2][2] ));
   NOR2 \mult_19_3/AN1_2_1  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[2][1] ));
   NOR2 \mult_19_3/AN1_2_0_0  (.A(\mult_19_3/A_notx [2]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[2][0] ));
   NOR2 \mult_19_3/AN2_1_7  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[1][7] ));
   NOR2 \mult_19_3/AN1_1_6  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[1][6] ));
   NOR2 \mult_19_3/AN1_1_5  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[1][5] ));
   NOR2 \mult_19_3/AN1_1_4  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[1][4] ));
   NOR2 \mult_19_3/AN1_1_3  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[1][3] ));
   NOR2 \mult_19_3/AN1_1_2  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[1][2] ));
   NOR2 \mult_19_3/AN1_1_1  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[1][1] ));
   NOR2 \mult_19_3/AN1_1_0_0  (.A(\mult_19_3/A_notx [1]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(\mult_19_3/ab[1][0] ));
   NOR2 \mult_19_3/AN2_0_7  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_not[7] ),
	.OUT(\mult_19_3/ab[0][7] ));
   NOR2 \mult_19_3/AN1_0_6  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [6]),
	.OUT(\mult_19_3/ab[0][6] ));
   NOR2 \mult_19_3/AN1_0_5  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [5]),
	.OUT(\mult_19_3/ab[0][5] ));
   NOR2 \mult_19_3/AN1_0_4  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [4]),
	.OUT(\mult_19_3/ab[0][4] ));
   NOR2 \mult_19_3/AN1_0_3  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [3]),
	.OUT(\mult_19_3/ab[0][3] ));
   NOR2 \mult_19_3/AN1_0_2  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [2]),
	.OUT(\mult_19_3/ab[0][2] ));
   NOR2 \mult_19_3/AN1_0_1  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [1]),
	.OUT(\mult_19_3/ab[0][1] ));
   NOR2 \mult_19_3/AN1_0_0_0  (.A(\mult_19_3/A_notx [0]),
	.B(\mult_19_3/B_notx [0]),
	.OUT(N49));
   OAI21 \mult_19_2/FS_1/U6_1_0_3  (.OUT(\mult_19_2/FS_1/C[1][3][0] ),
	.C(n2979),
	.B(n2978),
	.A(n2977));
   OAI21 \mult_19_2/FS_1/U6_0_3_1  (.OUT(\mult_19_2/FS_1/C[1][3][1] ),
	.C(\mult_19_2/FS_1/G_n_int[0][3][0] ),
	.B(n2975),
	.A(n2974));
   XOR2 \mult_19_2/FS_1/U3_C_0_3_1  (.A(\mult_19_2/FS_1/PG_int[0][3][1] ),
	.B(\mult_19_2/FS_1/C[1][3][1] ),
	.OUT(N32));
   XOR2 \mult_19_2/FS_1/U3_C_0_3_0  (.A(\mult_19_2/FS_1/PG_int[0][3][0] ),
	.B(\mult_19_2/FS_1/C[1][3][0] ),
	.OUT(N31));
   NAND2 \mult_19_2/FS_1/U3_B_0_3_0  (.A(\mult_19_2/FS_1/G_n_int[0][3][0] ),
	.B(\mult_19_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2971));
   NAND2 \mult_19_2/FS_1/U2_0_3_0  (.A(\mult_19_2/A1[12] ),
	.B(\mult_19_2/A2[12] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_19_2/FS_1/U1_0_3_0  (.A(n2969),
	.B(n2970),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_19_2/FS_1/U6_0_2_3  (.OUT(\mult_19_2/FS_1/C[1][2][3] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][2] ),
	.B(n2968),
	.A(n2967));
   OAI21 \mult_19_2/FS_1/U5_0_2_3  (.OUT(\mult_19_2/FS_1/G[1][0][2] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][3] ),
	.B(n2966),
	.A(n2965));
   NAND2 \mult_19_2/FS_1/U4_0_2_3  (.A(\mult_19_2/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_19_2/FS_1/P[0][2][3] ),
	.OUT(n2978));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_3  (.A(\mult_19_2/FS_1/PG_int[0][2][3] ),
	.B(\mult_19_2/FS_1/C[1][2][3] ),
	.OUT(N30));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_3  (.A(\mult_19_2/FS_1/G_n_int[0][2][3] ),
	.B(\mult_19_2/FS_1/P[0][2][3] ),
	.OUT(n2964));
   NAND2 \mult_19_2/FS_1/U2_0_2_3  (.A(\mult_19_2/A1[11] ),
	.B(\mult_19_2/A2[11] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_3  (.A(n2962),
	.B(n2963),
	.OUT(\mult_19_2/FS_1/P[0][2][3] ));
   OAI21 \mult_19_2/FS_1/U6_0_2_2  (.OUT(\mult_19_2/FS_1/C[1][2][2] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][1] ),
	.B(n2961),
	.A(n2960));
   OAI21 \mult_19_2/FS_1/U5_0_2_2  (.OUT(\mult_19_2/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][2] ),
	.B(n2968),
	.A(n2959));
   NAND2 \mult_19_2/FS_1/U4_0_2_2  (.A(\mult_19_2/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_19_2/FS_1/P[0][2][2] ),
	.OUT(n2958));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_2  (.A(\mult_19_2/FS_1/PG_int[0][2][2] ),
	.B(\mult_19_2/FS_1/C[1][2][2] ),
	.OUT(N29));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_2  (.A(\mult_19_2/FS_1/G_n_int[0][2][2] ),
	.B(\mult_19_2/FS_1/P[0][2][2] ),
	.OUT(n2957));
   NAND2 \mult_19_2/FS_1/U2_0_2_2  (.A(\mult_19_2/A1[10] ),
	.B(\mult_19_2/A2[10] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_2  (.A(n2955),
	.B(n2956),
	.OUT(\mult_19_2/FS_1/P[0][2][2] ));
   OAI21 \mult_19_2/FS_1/U6_0_2_1  (.OUT(\mult_19_2/FS_1/C[1][2][1] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][0] ),
	.B(n2954),
	.A(n2977));
   OAI21 \mult_19_2/FS_1/U5_0_2_1  (.OUT(\mult_19_2/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_19_2/FS_1/G_n_int[0][2][1] ),
	.B(n2961),
	.A(\mult_19_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_2/FS_1/U4_0_2_1  (.A(\mult_19_2/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_19_2/FS_1/P[0][2][1] ),
	.OUT(n2953));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_1  (.A(\mult_19_2/FS_1/PG_int[0][2][1] ),
	.B(\mult_19_2/FS_1/C[1][2][1] ),
	.OUT(N28));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_1  (.A(\mult_19_2/FS_1/G_n_int[0][2][1] ),
	.B(\mult_19_2/FS_1/P[0][2][1] ),
	.OUT(n2952));
   NAND2 \mult_19_2/FS_1/U2_0_2_1  (.A(\mult_19_2/A1[9] ),
	.B(\mult_19_2/A2[9] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_1  (.A(n2950),
	.B(n2951),
	.OUT(\mult_19_2/FS_1/P[0][2][1] ));
   XOR2 \mult_19_2/FS_1/U3_C_0_2_0  (.A(\mult_19_2/FS_1/PG_int[0][2][0] ),
	.B(\mult_19_2/FS_1/C[1][2][0] ),
	.OUT(N27));
   NAND2 \mult_19_2/FS_1/U3_B_0_2_0  (.A(\mult_19_2/FS_1/G_n_int[0][2][0] ),
	.B(\mult_19_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2949));
   NAND2 \mult_19_2/FS_1/U2_0_2_0  (.A(\mult_19_2/A1[8] ),
	.B(\mult_19_2/A2[8] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19_2/FS_1/U1_0_2_0  (.A(n2947),
	.B(n2948),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_19_2/FS_1/U3_B_0_1_3  (.A(\mult_19_2/FS_1/G_n_int[0][1][3] ),
	.B(\mult_19_2/FS_1/P[0][1][3] ),
	.OUT(n2946));
   NAND2 \mult_19_2/FS_1/U2_0_1_3  (.A(\mult_19_2/A1[7] ),
	.B(\mult_19_2/A2[7] ),
	.OUT(\mult_19_2/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_19_2/FS_1/U1_0_1_3  (.A(n2944),
	.B(n2945),
	.OUT(\mult_19_2/FS_1/P[0][1][3] ));
   INVERTER \mult_19_2/AN1_7  (.IN(matrix01[7]),
	.OUT(\mult_19_2/A_not[7] ));
   INVERTER \mult_19_2/AN1_6  (.IN(matrix01[6]),
	.OUT(\mult_19_2/A_notx [6]));
   INVERTER \mult_19_2/AN1_5  (.IN(matrix01[5]),
	.OUT(\mult_19_2/A_notx [5]));
   INVERTER \mult_19_2/AN1_4  (.IN(matrix01[4]),
	.OUT(\mult_19_2/A_notx [4]));
   INVERTER \mult_19_2/AN1_3  (.IN(matrix01[3]),
	.OUT(\mult_19_2/A_notx [3]));
   INVERTER \mult_19_2/AN1_2  (.IN(matrix01[2]),
	.OUT(\mult_19_2/A_notx [2]));
   INVERTER \mult_19_2/AN1_1  (.IN(matrix01[1]),
	.OUT(\mult_19_2/A_notx [1]));
   INVERTER \mult_19_2/AN1_0  (.IN(matrix01[0]),
	.OUT(\mult_19_2/A_notx [0]));
   INVERTER \mult_19_2/AN1_7_0  (.IN(vector_1[7]),
	.OUT(\mult_19_2/B_not[7] ));
   INVERTER \mult_19_2/AN1_6_0  (.IN(vector_1[6]),
	.OUT(\mult_19_2/B_notx [6]));
   INVERTER \mult_19_2/AN1_5_0  (.IN(vector_1[5]),
	.OUT(\mult_19_2/B_notx [5]));
   INVERTER \mult_19_2/AN1_4_0  (.IN(vector_1[4]),
	.OUT(\mult_19_2/B_notx [4]));
   INVERTER \mult_19_2/AN1_3_0  (.IN(vector_1[3]),
	.OUT(\mult_19_2/B_notx [3]));
   INVERTER \mult_19_2/AN1_2_0  (.IN(vector_1[2]),
	.OUT(\mult_19_2/B_notx [2]));
   INVERTER \mult_19_2/AN1_1_0  (.IN(vector_1[1]),
	.OUT(\mult_19_2/B_notx [1]));
   INVERTER \mult_19_2/AN1_0_0  (.IN(vector_1[0]),
	.OUT(\mult_19_2/B_notx [0]));
   NOR2 \mult_19_2/AN1_7_7  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[7][7] ));
   NOR2 \mult_19_2/AN3_7_6  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[7][6] ));
   NOR2 \mult_19_2/AN3_7_5  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[7][5] ));
   NOR2 \mult_19_2/AN3_7_4  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[7][4] ));
   NOR2 \mult_19_2/AN3_7_3  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[7][3] ));
   NOR2 \mult_19_2/AN3_7_2  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[7][2] ));
   NOR2 \mult_19_2/AN3_7_1  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[7][1] ));
   NOR2 \mult_19_2/AN3_7_0  (.A(\mult_19_2/A_not[7] ),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[7][0] ));
   NOR2 \mult_19_2/AN2_6_7  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[6][7] ));
   NOR2 \mult_19_2/AN1_6_6  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[6][6] ));
   NOR2 \mult_19_2/AN1_6_5  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[6][5] ));
   NOR2 \mult_19_2/AN1_6_4  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[6][4] ));
   NOR2 \mult_19_2/AN1_6_3  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[6][3] ));
   NOR2 \mult_19_2/AN1_6_2  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[6][2] ));
   NOR2 \mult_19_2/AN1_6_1  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[6][1] ));
   NOR2 \mult_19_2/AN1_6_0_0  (.A(\mult_19_2/A_notx [6]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[6][0] ));
   NOR2 \mult_19_2/AN2_5_7  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[5][7] ));
   NOR2 \mult_19_2/AN1_5_6  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[5][6] ));
   NOR2 \mult_19_2/AN1_5_5  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[5][5] ));
   NOR2 \mult_19_2/AN1_5_4  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[5][4] ));
   NOR2 \mult_19_2/AN1_5_3  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[5][3] ));
   NOR2 \mult_19_2/AN1_5_2  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[5][2] ));
   NOR2 \mult_19_2/AN1_5_1  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[5][1] ));
   NOR2 \mult_19_2/AN1_5_0_0  (.A(\mult_19_2/A_notx [5]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[5][0] ));
   NOR2 \mult_19_2/AN2_4_7  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[4][7] ));
   NOR2 \mult_19_2/AN1_4_6  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[4][6] ));
   NOR2 \mult_19_2/AN1_4_5  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[4][5] ));
   NOR2 \mult_19_2/AN1_4_4  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[4][4] ));
   NOR2 \mult_19_2/AN1_4_3  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[4][3] ));
   NOR2 \mult_19_2/AN1_4_2  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[4][2] ));
   NOR2 \mult_19_2/AN1_4_1  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[4][1] ));
   NOR2 \mult_19_2/AN1_4_0_0  (.A(\mult_19_2/A_notx [4]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[4][0] ));
   NOR2 \mult_19_2/AN2_3_7  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[3][7] ));
   NOR2 \mult_19_2/AN1_3_6  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[3][6] ));
   NOR2 \mult_19_2/AN1_3_5  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[3][5] ));
   NOR2 \mult_19_2/AN1_3_4  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[3][4] ));
   NOR2 \mult_19_2/AN1_3_3  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[3][3] ));
   NOR2 \mult_19_2/AN1_3_2  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[3][2] ));
   NOR2 \mult_19_2/AN1_3_1  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[3][1] ));
   NOR2 \mult_19_2/AN1_3_0_0  (.A(\mult_19_2/A_notx [3]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[3][0] ));
   NOR2 \mult_19_2/AN2_2_7  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[2][7] ));
   NOR2 \mult_19_2/AN1_2_6  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[2][6] ));
   NOR2 \mult_19_2/AN1_2_5  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[2][5] ));
   NOR2 \mult_19_2/AN1_2_4  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[2][4] ));
   NOR2 \mult_19_2/AN1_2_3  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[2][3] ));
   NOR2 \mult_19_2/AN1_2_2  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[2][2] ));
   NOR2 \mult_19_2/AN1_2_1  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[2][1] ));
   NOR2 \mult_19_2/AN1_2_0_0  (.A(\mult_19_2/A_notx [2]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[2][0] ));
   NOR2 \mult_19_2/AN2_1_7  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[1][7] ));
   NOR2 \mult_19_2/AN1_1_6  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[1][6] ));
   NOR2 \mult_19_2/AN1_1_5  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[1][5] ));
   NOR2 \mult_19_2/AN1_1_4  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[1][4] ));
   NOR2 \mult_19_2/AN1_1_3  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[1][3] ));
   NOR2 \mult_19_2/AN1_1_2  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[1][2] ));
   NOR2 \mult_19_2/AN1_1_1  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[1][1] ));
   NOR2 \mult_19_2/AN1_1_0_0  (.A(\mult_19_2/A_notx [1]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(\mult_19_2/ab[1][0] ));
   NOR2 \mult_19_2/AN2_0_7  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_not[7] ),
	.OUT(\mult_19_2/ab[0][7] ));
   NOR2 \mult_19_2/AN1_0_6  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [6]),
	.OUT(\mult_19_2/ab[0][6] ));
   NOR2 \mult_19_2/AN1_0_5  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [5]),
	.OUT(\mult_19_2/ab[0][5] ));
   NOR2 \mult_19_2/AN1_0_4  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [4]),
	.OUT(\mult_19_2/ab[0][4] ));
   NOR2 \mult_19_2/AN1_0_3  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [3]),
	.OUT(\mult_19_2/ab[0][3] ));
   NOR2 \mult_19_2/AN1_0_2  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [2]),
	.OUT(\mult_19_2/ab[0][2] ));
   NOR2 \mult_19_2/AN1_0_1  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [1]),
	.OUT(\mult_19_2/ab[0][1] ));
   NOR2 \mult_19_2/AN1_0_0_0  (.A(\mult_19_2/A_notx [0]),
	.B(\mult_19_2/B_notx [0]),
	.OUT(N17));
   OAI21 \mult_19/FS_1/U6_1_0_3  (.OUT(\mult_19/FS_1/C[1][3][0] ),
	.C(n2929),
	.B(n2928),
	.A(n2927));
   OAI21 \mult_19/FS_1/U6_0_3_1  (.OUT(\mult_19/FS_1/C[1][3][1] ),
	.C(\mult_19/FS_1/G_n_int[0][3][0] ),
	.B(n2925),
	.A(n2924));
   XOR2 \mult_19/FS_1/U3_C_0_3_1  (.A(\mult_19/FS_1/PG_int[0][3][1] ),
	.B(\mult_19/FS_1/C[1][3][1] ),
	.OUT(N16));
   XOR2 \mult_19/FS_1/U3_C_0_3_0  (.A(\mult_19/FS_1/PG_int[0][3][0] ),
	.B(\mult_19/FS_1/C[1][3][0] ),
	.OUT(N15));
   NAND2 \mult_19/FS_1/U3_B_0_3_0  (.A(\mult_19/FS_1/G_n_int[0][3][0] ),
	.B(\mult_19/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2921));
   NAND2 \mult_19/FS_1/U2_0_3_0  (.A(\mult_19/A1[12] ),
	.B(\mult_19/A2[12] ),
	.OUT(\mult_19/FS_1/G_n_int[0][3][0] ));
   NAND2 \mult_19/FS_1/U1_0_3_0  (.A(n2919),
	.B(n2920),
	.OUT(\mult_19/FS_1/TEMP_P[0][3][0] ));
   OAI21 \mult_19/FS_1/U6_0_2_3  (.OUT(\mult_19/FS_1/C[1][2][3] ),
	.C(\mult_19/FS_1/G_n_int[0][2][2] ),
	.B(n2918),
	.A(n2917));
   OAI21 \mult_19/FS_1/U5_0_2_3  (.OUT(\mult_19/FS_1/G[1][0][2] ),
	.C(\mult_19/FS_1/G_n_int[0][2][3] ),
	.B(n2916),
	.A(n2915));
   NAND2 \mult_19/FS_1/U4_0_2_3  (.A(\mult_19/FS_1/TEMP_P[0][2][2] ),
	.B(\mult_19/FS_1/P[0][2][3] ),
	.OUT(n2928));
   XOR2 \mult_19/FS_1/U3_C_0_2_3  (.A(\mult_19/FS_1/PG_int[0][2][3] ),
	.B(\mult_19/FS_1/C[1][2][3] ),
	.OUT(N14));
   NAND2 \mult_19/FS_1/U3_B_0_2_3  (.A(\mult_19/FS_1/G_n_int[0][2][3] ),
	.B(\mult_19/FS_1/P[0][2][3] ),
	.OUT(n2914));
   NAND2 \mult_19/FS_1/U2_0_2_3  (.A(\mult_19/A1[11] ),
	.B(\mult_19/A2[11] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][3] ));
   NAND2 \mult_19/FS_1/U1_0_2_3  (.A(n2912),
	.B(n2913),
	.OUT(\mult_19/FS_1/P[0][2][3] ));
   OAI21 \mult_19/FS_1/U6_0_2_2  (.OUT(\mult_19/FS_1/C[1][2][2] ),
	.C(\mult_19/FS_1/G_n_int[0][2][1] ),
	.B(n2911),
	.A(n2910));
   OAI21 \mult_19/FS_1/U5_0_2_2  (.OUT(\mult_19/FS_1/TEMP_G[0][2][2] ),
	.C(\mult_19/FS_1/G_n_int[0][2][2] ),
	.B(n2918),
	.A(n2909));
   NAND2 \mult_19/FS_1/U4_0_2_2  (.A(\mult_19/FS_1/TEMP_P[0][2][1] ),
	.B(\mult_19/FS_1/P[0][2][2] ),
	.OUT(n2908));
   XOR2 \mult_19/FS_1/U3_C_0_2_2  (.A(\mult_19/FS_1/PG_int[0][2][2] ),
	.B(\mult_19/FS_1/C[1][2][2] ),
	.OUT(N13));
   NAND2 \mult_19/FS_1/U3_B_0_2_2  (.A(\mult_19/FS_1/G_n_int[0][2][2] ),
	.B(\mult_19/FS_1/P[0][2][2] ),
	.OUT(n2907));
   NAND2 \mult_19/FS_1/U2_0_2_2  (.A(\mult_19/A1[10] ),
	.B(\mult_19/A2[10] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][2] ));
   NAND2 \mult_19/FS_1/U1_0_2_2  (.A(n2905),
	.B(n2906),
	.OUT(\mult_19/FS_1/P[0][2][2] ));
   OAI21 \mult_19/FS_1/U6_0_2_1  (.OUT(\mult_19/FS_1/C[1][2][1] ),
	.C(\mult_19/FS_1/G_n_int[0][2][0] ),
	.B(n2904),
	.A(n2927));
   OAI21 \mult_19/FS_1/U5_0_2_1  (.OUT(\mult_19/FS_1/TEMP_G[0][2][1] ),
	.C(\mult_19/FS_1/G_n_int[0][2][1] ),
	.B(n2911),
	.A(\mult_19/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19/FS_1/U4_0_2_1  (.A(\mult_19/FS_1/TEMP_P[0][2][0] ),
	.B(\mult_19/FS_1/P[0][2][1] ),
	.OUT(n2903));
   XOR2 \mult_19/FS_1/U3_C_0_2_1  (.A(\mult_19/FS_1/PG_int[0][2][1] ),
	.B(\mult_19/FS_1/C[1][2][1] ),
	.OUT(N12));
   NAND2 \mult_19/FS_1/U3_B_0_2_1  (.A(\mult_19/FS_1/G_n_int[0][2][1] ),
	.B(\mult_19/FS_1/P[0][2][1] ),
	.OUT(n2902));
   NAND2 \mult_19/FS_1/U2_0_2_1  (.A(\mult_19/A1[9] ),
	.B(\mult_19/A2[9] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][1] ));
   NAND2 \mult_19/FS_1/U1_0_2_1  (.A(n2900),
	.B(n2901),
	.OUT(\mult_19/FS_1/P[0][2][1] ));
   XOR2 \mult_19/FS_1/U3_C_0_2_0  (.A(\mult_19/FS_1/PG_int[0][2][0] ),
	.B(\mult_19/FS_1/C[1][2][0] ),
	.OUT(N11));
   NAND2 \mult_19/FS_1/U3_B_0_2_0  (.A(\mult_19/FS_1/G_n_int[0][2][0] ),
	.B(\mult_19/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2899));
   NAND2 \mult_19/FS_1/U2_0_2_0  (.A(\mult_19/A1[8] ),
	.B(\mult_19/A2[8] ),
	.OUT(\mult_19/FS_1/G_n_int[0][2][0] ));
   NAND2 \mult_19/FS_1/U1_0_2_0  (.A(n2897),
	.B(n2898),
	.OUT(\mult_19/FS_1/TEMP_P[0][2][0] ));
   NAND2 \mult_19/FS_1/U3_B_0_1_3  (.A(\mult_19/FS_1/G_n_int[0][1][3] ),
	.B(\mult_19/FS_1/P[0][1][3] ),
	.OUT(n2896));
   NAND2 \mult_19/FS_1/U2_0_1_3  (.A(\mult_19/A1[7] ),
	.B(\mult_19/A2[7] ),
	.OUT(\mult_19/FS_1/G_n_int[0][1][3] ));
   NAND2 \mult_19/FS_1/U1_0_1_3  (.A(n2894),
	.B(n2895),
	.OUT(\mult_19/FS_1/P[0][1][3] ));
   INVERTER \mult_19/AN1_7  (.IN(matrix00[7]),
	.OUT(\mult_19/A_not[7] ));
   INVERTER \mult_19/AN1_6  (.IN(matrix00[6]),
	.OUT(\mult_19/A_notx [6]));
   INVERTER \mult_19/AN1_5  (.IN(matrix00[5]),
	.OUT(\mult_19/A_notx [5]));
   INVERTER \mult_19/AN1_4  (.IN(matrix00[4]),
	.OUT(\mult_19/A_notx [4]));
   INVERTER \mult_19/AN1_3  (.IN(matrix00[3]),
	.OUT(\mult_19/A_notx [3]));
   INVERTER \mult_19/AN1_2  (.IN(matrix00[2]),
	.OUT(\mult_19/A_notx [2]));
   INVERTER \mult_19/AN1_1  (.IN(matrix00[1]),
	.OUT(\mult_19/A_notx [1]));
   INVERTER \mult_19/AN1_0  (.IN(matrix00[0]),
	.OUT(\mult_19/A_notx [0]));
   INVERTER \mult_19/AN1_7_0  (.IN(vector_0[7]),
	.OUT(\mult_19/B_not[7] ));
   INVERTER \mult_19/AN1_6_0  (.IN(vector_0[6]),
	.OUT(\mult_19/B_notx [6]));
   INVERTER \mult_19/AN1_5_0  (.IN(vector_0[5]),
	.OUT(\mult_19/B_notx [5]));
   INVERTER \mult_19/AN1_4_0  (.IN(vector_0[4]),
	.OUT(\mult_19/B_notx [4]));
   INVERTER \mult_19/AN1_3_0  (.IN(vector_0[3]),
	.OUT(\mult_19/B_notx [3]));
   INVERTER \mult_19/AN1_2_0  (.IN(vector_0[2]),
	.OUT(\mult_19/B_notx [2]));
   INVERTER \mult_19/AN1_1_0  (.IN(vector_0[1]),
	.OUT(\mult_19/B_notx [1]));
   INVERTER \mult_19/AN1_0_0  (.IN(vector_0[0]),
	.OUT(\mult_19/B_notx [0]));
   NOR2 \mult_19/AN1_7_7  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[7][7] ));
   NOR2 \mult_19/AN3_7_6  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[7][6] ));
   NOR2 \mult_19/AN3_7_5  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[7][5] ));
   NOR2 \mult_19/AN3_7_4  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[7][4] ));
   NOR2 \mult_19/AN3_7_3  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[7][3] ));
   NOR2 \mult_19/AN3_7_2  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[7][2] ));
   NOR2 \mult_19/AN3_7_1  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[7][1] ));
   NOR2 \mult_19/AN3_7_0  (.A(\mult_19/A_not[7] ),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[7][0] ));
   NOR2 \mult_19/AN2_6_7  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[6][7] ));
   NOR2 \mult_19/AN1_6_6  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[6][6] ));
   NOR2 \mult_19/AN1_6_5  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[6][5] ));
   NOR2 \mult_19/AN1_6_4  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[6][4] ));
   NOR2 \mult_19/AN1_6_3  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[6][3] ));
   NOR2 \mult_19/AN1_6_2  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[6][2] ));
   NOR2 \mult_19/AN1_6_1  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[6][1] ));
   NOR2 \mult_19/AN1_6_0_0  (.A(\mult_19/A_notx [6]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[6][0] ));
   NOR2 \mult_19/AN2_5_7  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[5][7] ));
   NOR2 \mult_19/AN1_5_6  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[5][6] ));
   NOR2 \mult_19/AN1_5_5  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[5][5] ));
   NOR2 \mult_19/AN1_5_4  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[5][4] ));
   NOR2 \mult_19/AN1_5_3  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[5][3] ));
   NOR2 \mult_19/AN1_5_2  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[5][2] ));
   NOR2 \mult_19/AN1_5_1  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[5][1] ));
   NOR2 \mult_19/AN1_5_0_0  (.A(\mult_19/A_notx [5]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[5][0] ));
   NOR2 \mult_19/AN2_4_7  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[4][7] ));
   NOR2 \mult_19/AN1_4_6  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[4][6] ));
   NOR2 \mult_19/AN1_4_5  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[4][5] ));
   NOR2 \mult_19/AN1_4_4  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[4][4] ));
   NOR2 \mult_19/AN1_4_3  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[4][3] ));
   NOR2 \mult_19/AN1_4_2  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[4][2] ));
   NOR2 \mult_19/AN1_4_1  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[4][1] ));
   NOR2 \mult_19/AN1_4_0_0  (.A(\mult_19/A_notx [4]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[4][0] ));
   NOR2 \mult_19/AN2_3_7  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[3][7] ));
   NOR2 \mult_19/AN1_3_6  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[3][6] ));
   NOR2 \mult_19/AN1_3_5  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[3][5] ));
   NOR2 \mult_19/AN1_3_4  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[3][4] ));
   NOR2 \mult_19/AN1_3_3  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[3][3] ));
   NOR2 \mult_19/AN1_3_2  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[3][2] ));
   NOR2 \mult_19/AN1_3_1  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[3][1] ));
   NOR2 \mult_19/AN1_3_0_0  (.A(\mult_19/A_notx [3]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[3][0] ));
   NOR2 \mult_19/AN2_2_7  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[2][7] ));
   NOR2 \mult_19/AN1_2_6  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[2][6] ));
   NOR2 \mult_19/AN1_2_5  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[2][5] ));
   NOR2 \mult_19/AN1_2_4  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[2][4] ));
   NOR2 \mult_19/AN1_2_3  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[2][3] ));
   NOR2 \mult_19/AN1_2_2  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[2][2] ));
   NOR2 \mult_19/AN1_2_1  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[2][1] ));
   NOR2 \mult_19/AN1_2_0_0  (.A(\mult_19/A_notx [2]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[2][0] ));
   NOR2 \mult_19/AN2_1_7  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[1][7] ));
   NOR2 \mult_19/AN1_1_6  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[1][6] ));
   NOR2 \mult_19/AN1_1_5  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[1][5] ));
   NOR2 \mult_19/AN1_1_4  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[1][4] ));
   NOR2 \mult_19/AN1_1_3  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[1][3] ));
   NOR2 \mult_19/AN1_1_2  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[1][2] ));
   NOR2 \mult_19/AN1_1_1  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[1][1] ));
   NOR2 \mult_19/AN1_1_0_0  (.A(\mult_19/A_notx [1]),
	.B(\mult_19/B_notx [0]),
	.OUT(\mult_19/ab[1][0] ));
   NOR2 \mult_19/AN2_0_7  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_not[7] ),
	.OUT(\mult_19/ab[0][7] ));
   NOR2 \mult_19/AN1_0_6  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [6]),
	.OUT(\mult_19/ab[0][6] ));
   NOR2 \mult_19/AN1_0_5  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [5]),
	.OUT(\mult_19/ab[0][5] ));
   NOR2 \mult_19/AN1_0_4  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [4]),
	.OUT(\mult_19/ab[0][4] ));
   NOR2 \mult_19/AN1_0_3  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [3]),
	.OUT(\mult_19/ab[0][3] ));
   NOR2 \mult_19/AN1_0_2  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [2]),
	.OUT(\mult_19/ab[0][2] ));
   NOR2 \mult_19/AN1_0_1  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [1]),
	.OUT(\mult_19/ab[0][1] ));
   NOR2 \mult_19/AN1_0_0_0  (.A(\mult_19/A_notx [0]),
	.B(\mult_19/B_notx [0]),
	.OUT(N1));
   INVERTER U19 (.IN(clk),
	.OUT(n17));
   INVERTER U20 (.IN(clk),
	.OUT(n18));
   INVERTER U21 (.IN(clk),
	.OUT(n19));
   INVERTER U22 (.IN(clk),
	.OUT(n20));
   INVERTER U23 (.IN(clk),
	.OUT(n21));
   INVERTER U24 (.IN(clk),
	.OUT(n22));
   INVERTER U25 (.IN(clk),
	.OUT(n23));
   INVERTER U26 (.IN(clk),
	.OUT(n24));
   INVERTER U27 (.IN(clk),
	.OUT(n25));
   INVERTER U28 (.IN(clk),
	.OUT(n26));
   INVERTER U29 (.IN(clk),
	.OUT(n27));
   INVERTER U30 (.IN(clk),
	.OUT(n28));
   INVERTER U31 (.IN(clk),
	.OUT(n29));
   INVERTER U32 (.IN(clk),
	.OUT(n30));
   INVERTER U33 (.IN(clk),
	.OUT(n31));
   INVERTER U34 (.IN(clk),
	.OUT(n32));
   INVERTER U35 (.IN(clk),
	.OUT(n33));
   INVERTER U36 (.IN(clk),
	.OUT(n34));
   INVERTER U37 (.IN(clk),
	.OUT(n35));
   INVERTER U38 (.IN(clk),
	.OUT(n36));
   INVERTER U39 (.IN(clk),
	.OUT(n37));
   INVERTER U40 (.IN(clk),
	.OUT(n38));
   INVERTER U41 (.IN(clk),
	.OUT(n39));
   INVERTER U42 (.IN(clk),
	.OUT(n40));
   INVERTER U43 (.IN(clk),
	.OUT(n41));
   INVERTER U44 (.IN(clk),
	.OUT(n42));
   INVERTER U45 (.IN(clk),
	.OUT(n43));
   INVERTER U46 (.IN(clk),
	.OUT(n44));
   INVERTER U47 (.IN(clk),
	.OUT(n45));
   INVERTER U48 (.IN(clk),
	.OUT(n46));
   INVERTER U49 (.IN(clk),
	.OUT(n47));
   INVERTER U50 (.IN(clk),
	.OUT(n48));
   INVERTER U51 (.IN(clk),
	.OUT(n49));
   INVERTER U52 (.IN(clk),
	.OUT(n50));
   INVERTER U53 (.IN(clk),
	.OUT(n51));
   INVERTER U54 (.IN(clk),
	.OUT(n52));
   INVERTER U55 (.IN(clk),
	.OUT(n53));
   INVERTER U56 (.IN(rst_n),
	.OUT(n54));
   INVERTER U57 (.IN(rst_n),
	.OUT(n55));
   INVERTER U58 (.IN(clk),
	.OUT(n56));
   INVERTER U59 (.IN(clk),
	.OUT(n57));
   INVERTER U60 (.IN(clk),
	.OUT(n58));
   INVERTER U61 (.IN(clk),
	.OUT(n59));
   INVERTER U62 (.IN(clk),
	.OUT(n60));
   INVERTER U63 (.IN(clk),
	.OUT(n61));
   INVERTER U64 (.IN(clk),
	.OUT(n62));
   INVERTER U65 (.IN(clk),
	.OUT(n63));
   INVERTER U66 (.IN(clk),
	.OUT(n64));
   INVERTER U67 (.IN(clk),
	.OUT(n65));
   INVERTER U68 (.IN(n2880),
	.OUT(\mult_19/FS_1/TEMP_P[0][0][0] ));
   INVERTER U69 (.IN(n2930),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][0][0] ));
   INVERTER U70 (.IN(n2980),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][0][0] ));
   INVERTER U71 (.IN(n3030),
	.OUT(\mult_20/FS_1/TEMP_P[0][0][0] ));
   INVERTER U72 (.IN(n3080),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][0][0] ));
   INVERTER U73 (.IN(n3130),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][0][0] ));
   INVERTER U74 (.IN(n3180),
	.OUT(\mult_21/FS_1/TEMP_P[0][0][0] ));
   INVERTER U75 (.IN(n3230),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][0][0] ));
   INVERTER U76 (.IN(n3280),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][0][0] ));
   INVERTER U77 (.IN(\mult_21_3/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3281));
   INVERTER U78 (.IN(n3282),
	.OUT(\mult_21_3/FS_1/P[0][0][1] ));
   INVERTER U79 (.IN(\mult_21_3/FS_1/P[0][0][1] ),
	.OUT(n3283));
   INVERTER U80 (.IN(n3284),
	.OUT(\mult_21_3/FS_1/P[0][0][2] ));
   INVERTER U81 (.IN(\mult_21_3/FS_1/P[0][0][2] ),
	.OUT(n3285));
   INVERTER U82 (.IN(n3286),
	.OUT(\mult_21_3/FS_1/P[0][0][3] ));
   INVERTER U83 (.IN(\mult_21_3/FS_1/P[0][0][3] ),
	.OUT(n3287));
   INVERTER U84 (.IN(n3326),
	.OUT(\mult_21_3/FS_1/C[1][2][0] ));
   INVERTER U85 (.IN(n3288),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][1][0] ));
   INVERTER U86 (.IN(\mult_21_3/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3289));
   INVERTER U87 (.IN(n3290),
	.OUT(\mult_21_3/FS_1/P[0][1][1] ));
   INVERTER U88 (.IN(n3322),
	.OUT(\mult_21_3/FS_1/P[0][3][1] ));
   INVERTER U89 (.IN(\mult_21_3/FS_1/P[0][3][1] ),
	.OUT(n3323));
   INVERTER U90 (.IN(\mult_21_3/FS_1/P[0][1][1] ),
	.OUT(n3291));
   INVERTER U91 (.IN(n3292),
	.OUT(\mult_21_3/FS_1/P[0][1][2] ));
   INVERTER U92 (.IN(\mult_21_3/FS_1/P[0][1][2] ),
	.OUT(n3293));
   INVERTER U93 (.IN(\mult_21_3/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_21_3/FS_1/G[1][0][1] ));
   INVERTER U94 (.IN(\mult_21_2/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3231));
   INVERTER U95 (.IN(n3232),
	.OUT(\mult_21_2/FS_1/P[0][0][1] ));
   INVERTER U96 (.IN(\mult_21_2/FS_1/P[0][0][1] ),
	.OUT(n3233));
   INVERTER U97 (.IN(n3234),
	.OUT(\mult_21_2/FS_1/P[0][0][2] ));
   INVERTER U98 (.IN(\mult_21_2/FS_1/P[0][0][2] ),
	.OUT(n3235));
   INVERTER U99 (.IN(n3236),
	.OUT(\mult_21_2/FS_1/P[0][0][3] ));
   INVERTER U100 (.IN(\mult_21_2/FS_1/P[0][0][3] ),
	.OUT(n3237));
   INVERTER U101 (.IN(n3276),
	.OUT(\mult_21_2/FS_1/C[1][2][0] ));
   INVERTER U102 (.IN(n3238),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][1][0] ));
   INVERTER U103 (.IN(\mult_21_2/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3239));
   INVERTER U104 (.IN(n3240),
	.OUT(\mult_21_2/FS_1/P[0][1][1] ));
   INVERTER U105 (.IN(n3272),
	.OUT(\mult_21_2/FS_1/P[0][3][1] ));
   INVERTER U106 (.IN(\mult_21_2/FS_1/P[0][3][1] ),
	.OUT(n3273));
   INVERTER U107 (.IN(\mult_21_2/FS_1/P[0][1][1] ),
	.OUT(n3241));
   INVERTER U108 (.IN(n3242),
	.OUT(\mult_21_2/FS_1/P[0][1][2] ));
   INVERTER U109 (.IN(\mult_21_2/FS_1/P[0][1][2] ),
	.OUT(n3243));
   INVERTER U110 (.IN(\mult_21_2/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_21_2/FS_1/G[1][0][1] ));
   INVERTER U111 (.IN(\mult_21/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3181));
   INVERTER U112 (.IN(n3182),
	.OUT(\mult_21/FS_1/P[0][0][1] ));
   INVERTER U113 (.IN(\mult_21/FS_1/P[0][0][1] ),
	.OUT(n3183));
   INVERTER U114 (.IN(n3184),
	.OUT(\mult_21/FS_1/P[0][0][2] ));
   INVERTER U115 (.IN(\mult_21/FS_1/P[0][0][2] ),
	.OUT(n3185));
   INVERTER U116 (.IN(n3186),
	.OUT(\mult_21/FS_1/P[0][0][3] ));
   INVERTER U117 (.IN(\mult_21/FS_1/P[0][0][3] ),
	.OUT(n3187));
   INVERTER U118 (.IN(n3226),
	.OUT(\mult_21/FS_1/C[1][2][0] ));
   INVERTER U119 (.IN(n3188),
	.OUT(\mult_21/FS_1/TEMP_P[0][1][0] ));
   INVERTER U120 (.IN(\mult_21/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3189));
   INVERTER U121 (.IN(n3190),
	.OUT(\mult_21/FS_1/P[0][1][1] ));
   INVERTER U122 (.IN(n3222),
	.OUT(\mult_21/FS_1/P[0][3][1] ));
   INVERTER U123 (.IN(\mult_21/FS_1/P[0][3][1] ),
	.OUT(n3223));
   INVERTER U124 (.IN(\mult_21/FS_1/P[0][1][1] ),
	.OUT(n3191));
   INVERTER U125 (.IN(n3192),
	.OUT(\mult_21/FS_1/P[0][1][2] ));
   INVERTER U126 (.IN(\mult_21/FS_1/P[0][1][2] ),
	.OUT(n3193));
   INVERTER U127 (.IN(\mult_21/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_21/FS_1/G[1][0][1] ));
   INVERTER U128 (.IN(\mult_20_3/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3131));
   INVERTER U129 (.IN(n3132),
	.OUT(\mult_20_3/FS_1/P[0][0][1] ));
   INVERTER U130 (.IN(\mult_20_3/FS_1/P[0][0][1] ),
	.OUT(n3133));
   INVERTER U131 (.IN(n3134),
	.OUT(\mult_20_3/FS_1/P[0][0][2] ));
   INVERTER U132 (.IN(\mult_20_3/FS_1/P[0][0][2] ),
	.OUT(n3135));
   INVERTER U133 (.IN(n3136),
	.OUT(\mult_20_3/FS_1/P[0][0][3] ));
   INVERTER U134 (.IN(\mult_20_3/FS_1/P[0][0][3] ),
	.OUT(n3137));
   INVERTER U135 (.IN(n3176),
	.OUT(\mult_20_3/FS_1/C[1][2][0] ));
   INVERTER U136 (.IN(n3138),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][1][0] ));
   INVERTER U137 (.IN(\mult_20_3/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3139));
   INVERTER U138 (.IN(n3140),
	.OUT(\mult_20_3/FS_1/P[0][1][1] ));
   INVERTER U139 (.IN(n3172),
	.OUT(\mult_20_3/FS_1/P[0][3][1] ));
   INVERTER U140 (.IN(\mult_20_3/FS_1/P[0][3][1] ),
	.OUT(n3173));
   INVERTER U141 (.IN(\mult_20_3/FS_1/P[0][1][1] ),
	.OUT(n3141));
   INVERTER U142 (.IN(n3142),
	.OUT(\mult_20_3/FS_1/P[0][1][2] ));
   INVERTER U143 (.IN(\mult_20_3/FS_1/P[0][1][2] ),
	.OUT(n3143));
   INVERTER U144 (.IN(\mult_20_3/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_20_3/FS_1/G[1][0][1] ));
   INVERTER U145 (.IN(\mult_20_2/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3081));
   INVERTER U146 (.IN(n3082),
	.OUT(\mult_20_2/FS_1/P[0][0][1] ));
   INVERTER U147 (.IN(\mult_20_2/FS_1/P[0][0][1] ),
	.OUT(n3083));
   INVERTER U148 (.IN(n3084),
	.OUT(\mult_20_2/FS_1/P[0][0][2] ));
   INVERTER U149 (.IN(\mult_20_2/FS_1/P[0][0][2] ),
	.OUT(n3085));
   INVERTER U150 (.IN(n3086),
	.OUT(\mult_20_2/FS_1/P[0][0][3] ));
   INVERTER U151 (.IN(\mult_20_2/FS_1/P[0][0][3] ),
	.OUT(n3087));
   INVERTER U152 (.IN(n3126),
	.OUT(\mult_20_2/FS_1/C[1][2][0] ));
   INVERTER U153 (.IN(n3088),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][1][0] ));
   INVERTER U154 (.IN(\mult_20_2/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3089));
   INVERTER U155 (.IN(n3090),
	.OUT(\mult_20_2/FS_1/P[0][1][1] ));
   INVERTER U156 (.IN(n3122),
	.OUT(\mult_20_2/FS_1/P[0][3][1] ));
   INVERTER U157 (.IN(\mult_20_2/FS_1/P[0][3][1] ),
	.OUT(n3123));
   INVERTER U158 (.IN(\mult_20_2/FS_1/P[0][1][1] ),
	.OUT(n3091));
   INVERTER U159 (.IN(n3092),
	.OUT(\mult_20_2/FS_1/P[0][1][2] ));
   INVERTER U160 (.IN(\mult_20_2/FS_1/P[0][1][2] ),
	.OUT(n3093));
   INVERTER U161 (.IN(\mult_20_2/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_20_2/FS_1/G[1][0][1] ));
   INVERTER U162 (.IN(\mult_20/FS_1/TEMP_P[0][0][0] ),
	.OUT(n3031));
   INVERTER U163 (.IN(n3032),
	.OUT(\mult_20/FS_1/P[0][0][1] ));
   INVERTER U164 (.IN(\mult_20/FS_1/P[0][0][1] ),
	.OUT(n3033));
   INVERTER U165 (.IN(n3034),
	.OUT(\mult_20/FS_1/P[0][0][2] ));
   INVERTER U166 (.IN(\mult_20/FS_1/P[0][0][2] ),
	.OUT(n3035));
   INVERTER U167 (.IN(n3036),
	.OUT(\mult_20/FS_1/P[0][0][3] ));
   INVERTER U168 (.IN(\mult_20/FS_1/P[0][0][3] ),
	.OUT(n3037));
   INVERTER U169 (.IN(n3076),
	.OUT(\mult_20/FS_1/C[1][2][0] ));
   INVERTER U170 (.IN(n3038),
	.OUT(\mult_20/FS_1/TEMP_P[0][1][0] ));
   INVERTER U171 (.IN(\mult_20/FS_1/TEMP_P[0][1][0] ),
	.OUT(n3039));
   INVERTER U172 (.IN(n3040),
	.OUT(\mult_20/FS_1/P[0][1][1] ));
   INVERTER U173 (.IN(n3072),
	.OUT(\mult_20/FS_1/P[0][3][1] ));
   INVERTER U174 (.IN(\mult_20/FS_1/P[0][3][1] ),
	.OUT(n3073));
   INVERTER U175 (.IN(\mult_20/FS_1/P[0][1][1] ),
	.OUT(n3041));
   INVERTER U176 (.IN(n3042),
	.OUT(\mult_20/FS_1/P[0][1][2] ));
   INVERTER U177 (.IN(\mult_20/FS_1/P[0][1][2] ),
	.OUT(n3043));
   INVERTER U178 (.IN(\mult_20/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_20/FS_1/G[1][0][1] ));
   INVERTER U179 (.IN(\mult_19_3/FS_1/TEMP_P[0][0][0] ),
	.OUT(n2981));
   INVERTER U180 (.IN(n2982),
	.OUT(\mult_19_3/FS_1/P[0][0][1] ));
   INVERTER U181 (.IN(\mult_19_3/FS_1/P[0][0][1] ),
	.OUT(n2983));
   INVERTER U182 (.IN(n2984),
	.OUT(\mult_19_3/FS_1/P[0][0][2] ));
   INVERTER U183 (.IN(\mult_19_3/FS_1/P[0][0][2] ),
	.OUT(n2985));
   INVERTER U184 (.IN(n2986),
	.OUT(\mult_19_3/FS_1/P[0][0][3] ));
   INVERTER U185 (.IN(\mult_19_3/FS_1/P[0][0][3] ),
	.OUT(n2987));
   INVERTER U186 (.IN(n3026),
	.OUT(\mult_19_3/FS_1/C[1][2][0] ));
   INVERTER U187 (.IN(n2988),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][1][0] ));
   INVERTER U188 (.IN(\mult_19_3/FS_1/TEMP_P[0][1][0] ),
	.OUT(n2989));
   INVERTER U189 (.IN(n2990),
	.OUT(\mult_19_3/FS_1/P[0][1][1] ));
   INVERTER U190 (.IN(n3022),
	.OUT(\mult_19_3/FS_1/P[0][3][1] ));
   INVERTER U191 (.IN(\mult_19_3/FS_1/P[0][3][1] ),
	.OUT(n3023));
   INVERTER U192 (.IN(\mult_19_3/FS_1/P[0][1][1] ),
	.OUT(n2991));
   INVERTER U193 (.IN(n2992),
	.OUT(\mult_19_3/FS_1/P[0][1][2] ));
   INVERTER U194 (.IN(\mult_19_3/FS_1/P[0][1][2] ),
	.OUT(n2993));
   INVERTER U195 (.IN(\mult_19_3/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_19_3/FS_1/G[1][0][1] ));
   INVERTER U196 (.IN(\mult_19_2/FS_1/TEMP_P[0][0][0] ),
	.OUT(n2931));
   INVERTER U197 (.IN(n2932),
	.OUT(\mult_19_2/FS_1/P[0][0][1] ));
   INVERTER U198 (.IN(\mult_19_2/FS_1/P[0][0][1] ),
	.OUT(n2933));
   INVERTER U199 (.IN(n2934),
	.OUT(\mult_19_2/FS_1/P[0][0][2] ));
   INVERTER U200 (.IN(\mult_19_2/FS_1/P[0][0][2] ),
	.OUT(n2935));
   INVERTER U201 (.IN(n2936),
	.OUT(\mult_19_2/FS_1/P[0][0][3] ));
   INVERTER U202 (.IN(\mult_19_2/FS_1/P[0][0][3] ),
	.OUT(n2937));
   INVERTER U203 (.IN(n2976),
	.OUT(\mult_19_2/FS_1/C[1][2][0] ));
   INVERTER U204 (.IN(n2938),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][1][0] ));
   INVERTER U205 (.IN(\mult_19_2/FS_1/TEMP_P[0][1][0] ),
	.OUT(n2939));
   INVERTER U206 (.IN(n2940),
	.OUT(\mult_19_2/FS_1/P[0][1][1] ));
   INVERTER U207 (.IN(n2972),
	.OUT(\mult_19_2/FS_1/P[0][3][1] ));
   INVERTER U208 (.IN(\mult_19_2/FS_1/P[0][3][1] ),
	.OUT(n2973));
   INVERTER U209 (.IN(\mult_19_2/FS_1/P[0][1][1] ),
	.OUT(n2941));
   INVERTER U210 (.IN(n2942),
	.OUT(\mult_19_2/FS_1/P[0][1][2] ));
   INVERTER U211 (.IN(\mult_19_2/FS_1/P[0][1][2] ),
	.OUT(n2943));
   INVERTER U212 (.IN(\mult_19_2/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_19_2/FS_1/G[1][0][1] ));
   INVERTER U213 (.IN(\mult_19/FS_1/TEMP_P[0][0][0] ),
	.OUT(n2881));
   INVERTER U214 (.IN(n2882),
	.OUT(\mult_19/FS_1/P[0][0][1] ));
   INVERTER U215 (.IN(\mult_19/FS_1/P[0][0][1] ),
	.OUT(n2883));
   INVERTER U216 (.IN(n2884),
	.OUT(\mult_19/FS_1/P[0][0][2] ));
   INVERTER U217 (.IN(\mult_19/FS_1/P[0][0][2] ),
	.OUT(n2885));
   INVERTER U218 (.IN(n2886),
	.OUT(\mult_19/FS_1/P[0][0][3] ));
   INVERTER U219 (.IN(\mult_19/FS_1/P[0][0][3] ),
	.OUT(n2887));
   INVERTER U220 (.IN(n2926),
	.OUT(\mult_19/FS_1/C[1][2][0] ));
   INVERTER U221 (.IN(n2888),
	.OUT(\mult_19/FS_1/TEMP_P[0][1][0] ));
   INVERTER U222 (.IN(\mult_19/FS_1/TEMP_P[0][1][0] ),
	.OUT(n2889));
   INVERTER U223 (.IN(n2890),
	.OUT(\mult_19/FS_1/P[0][1][1] ));
   INVERTER U224 (.IN(n2922),
	.OUT(\mult_19/FS_1/P[0][3][1] ));
   INVERTER U225 (.IN(\mult_19/FS_1/P[0][3][1] ),
	.OUT(n2923));
   INVERTER U226 (.IN(\mult_19/FS_1/P[0][1][1] ),
	.OUT(n2891));
   INVERTER U227 (.IN(n2892),
	.OUT(\mult_19/FS_1/P[0][1][2] ));
   INVERTER U228 (.IN(\mult_19/FS_1/P[0][1][2] ),
	.OUT(n2893));
   INVERTER U229 (.IN(\mult_19/FS_1/G_n_int[0][1][3] ),
	.OUT(\mult_19/FS_1/G[1][0][1] ));
   NOR2 U230 (.A(n66),
	.B(n67),
	.OUT(\mult_19/A2[13] ));
   NAND2 U231 (.A(n69),
	.B(n70),
	.OUT(n68));
   NAND2 U232 (.A(n72),
	.B(n73),
	.OUT(n71));
   NOR2 U233 (.A(n74),
	.B(n75),
	.OUT(\mult_19/A2[10] ));
   NOR2 U234 (.A(n76),
	.B(n77),
	.OUT(\mult_19/A2[9] ));
   NOR2 U235 (.A(n78),
	.B(n79),
	.OUT(\mult_19/A2[8] ));
   NOR2 U236 (.A(n80),
	.B(n81),
	.OUT(\mult_19/A2[7] ));
   NOR2 U237 (.A(n82),
	.B(n83),
	.OUT(\mult_19_2/A2[13] ));
   NAND2 U238 (.A(n85),
	.B(n86),
	.OUT(n84));
   NAND2 U239 (.A(n88),
	.B(n89),
	.OUT(n87));
   NOR2 U240 (.A(n90),
	.B(n91),
	.OUT(\mult_19_2/A2[10] ));
   NOR2 U241 (.A(n92),
	.B(n93),
	.OUT(\mult_19_2/A2[9] ));
   NOR2 U242 (.A(n94),
	.B(n95),
	.OUT(\mult_19_2/A2[8] ));
   NOR2 U243 (.A(n96),
	.B(n97),
	.OUT(\mult_19_2/A2[7] ));
   NOR2 U244 (.A(n98),
	.B(n99),
	.OUT(\mult_19_3/A2[13] ));
   NAND2 U245 (.A(n101),
	.B(n102),
	.OUT(n100));
   NAND2 U246 (.A(n104),
	.B(n105),
	.OUT(n103));
   NOR2 U247 (.A(n106),
	.B(n107),
	.OUT(\mult_19_3/A2[10] ));
   NOR2 U248 (.A(n108),
	.B(n109),
	.OUT(\mult_19_3/A2[9] ));
   NOR2 U249 (.A(n110),
	.B(n111),
	.OUT(\mult_19_3/A2[8] ));
   NOR2 U250 (.A(n112),
	.B(n113),
	.OUT(\mult_19_3/A2[7] ));
   NOR2 U251 (.A(n114),
	.B(n115),
	.OUT(\mult_20/A2[13] ));
   NAND2 U252 (.A(n117),
	.B(n118),
	.OUT(n116));
   NAND2 U253 (.A(n120),
	.B(n121),
	.OUT(n119));
   NOR2 U254 (.A(n122),
	.B(n123),
	.OUT(\mult_20/A2[10] ));
   NOR2 U255 (.A(n124),
	.B(n125),
	.OUT(\mult_20/A2[9] ));
   NOR2 U256 (.A(n126),
	.B(n127),
	.OUT(\mult_20/A2[8] ));
   NOR2 U257 (.A(n128),
	.B(n129),
	.OUT(\mult_20/A2[7] ));
   NOR2 U258 (.A(n130),
	.B(n131),
	.OUT(\mult_20_2/A2[13] ));
   NAND2 U259 (.A(n133),
	.B(n134),
	.OUT(n132));
   NAND2 U260 (.A(n136),
	.B(n137),
	.OUT(n135));
   NOR2 U261 (.A(n138),
	.B(n139),
	.OUT(\mult_20_2/A2[10] ));
   NOR2 U262 (.A(n140),
	.B(n141),
	.OUT(\mult_20_2/A2[9] ));
   NOR2 U263 (.A(n142),
	.B(n143),
	.OUT(\mult_20_2/A2[8] ));
   NOR2 U264 (.A(n144),
	.B(n145),
	.OUT(\mult_20_2/A2[7] ));
   NOR2 U265 (.A(n146),
	.B(n147),
	.OUT(\mult_20_3/A2[13] ));
   NAND2 U266 (.A(n149),
	.B(n150),
	.OUT(n148));
   NAND2 U267 (.A(n152),
	.B(n153),
	.OUT(n151));
   NOR2 U268 (.A(n154),
	.B(n155),
	.OUT(\mult_20_3/A2[10] ));
   NOR2 U269 (.A(n156),
	.B(n157),
	.OUT(\mult_20_3/A2[9] ));
   NOR2 U270 (.A(n158),
	.B(n159),
	.OUT(\mult_20_3/A2[8] ));
   NOR2 U271 (.A(n160),
	.B(n161),
	.OUT(\mult_20_3/A2[7] ));
   NOR2 U272 (.A(n162),
	.B(n163),
	.OUT(\mult_21/A2[13] ));
   NAND2 U273 (.A(n165),
	.B(n166),
	.OUT(n164));
   NAND2 U274 (.A(n168),
	.B(n169),
	.OUT(n167));
   NOR2 U275 (.A(n170),
	.B(n171),
	.OUT(\mult_21/A2[10] ));
   NOR2 U276 (.A(n172),
	.B(n173),
	.OUT(\mult_21/A2[9] ));
   NOR2 U277 (.A(n174),
	.B(n175),
	.OUT(\mult_21/A2[8] ));
   NOR2 U278 (.A(n176),
	.B(n177),
	.OUT(\mult_21/A2[7] ));
   NOR2 U279 (.A(n178),
	.B(n179),
	.OUT(\mult_21_2/A2[13] ));
   NAND2 U280 (.A(n181),
	.B(n182),
	.OUT(n180));
   NAND2 U281 (.A(n184),
	.B(n185),
	.OUT(n183));
   NOR2 U282 (.A(n186),
	.B(n187),
	.OUT(\mult_21_2/A2[10] ));
   NOR2 U283 (.A(n188),
	.B(n189),
	.OUT(\mult_21_2/A2[9] ));
   NOR2 U284 (.A(n190),
	.B(n191),
	.OUT(\mult_21_2/A2[8] ));
   NOR2 U285 (.A(n192),
	.B(n193),
	.OUT(\mult_21_2/A2[7] ));
   NOR2 U286 (.A(n194),
	.B(n195),
	.OUT(\mult_21_3/A2[13] ));
   NAND2 U287 (.A(n197),
	.B(n198),
	.OUT(n196));
   NAND2 U288 (.A(n200),
	.B(n201),
	.OUT(n199));
   NOR2 U289 (.A(n202),
	.B(n203),
	.OUT(\mult_21_3/A2[10] ));
   NOR2 U290 (.A(n204),
	.B(n205),
	.OUT(\mult_21_3/A2[9] ));
   NOR2 U291 (.A(n206),
	.B(n207),
	.OUT(\mult_21_3/A2[8] ));
   NOR2 U292 (.A(n208),
	.B(n209),
	.OUT(\mult_21_3/A2[7] ));
   NOR2 U293 (.A(\mult_21_3/ab[1][7] ),
	.B(\mult_21_3/ab[2][6] ),
	.OUT(n210));
   NAND2 U294 (.A(n212),
	.B(n213),
	.OUT(n211));
   NOR2 U295 (.A(\mult_21_3/ab[4][5] ),
	.B(n215),
	.OUT(n214));
   NAND2 U296 (.A(n217),
	.B(n218),
	.OUT(n216));
   NOR2 U297 (.A(\mult_21_3/ab[4][4] ),
	.B(n220),
	.OUT(n219));
   NAND2 U298 (.A(n222),
	.B(n223),
	.OUT(n221));
   NOR2 U299 (.A(\mult_21_3/ab[4][3] ),
	.B(n225),
	.OUT(n224));
   NOR2 U300 (.A(\mult_21_3/ab[6][3] ),
	.B(n227),
	.OUT(n226));
   NOR2 U301 (.A(\mult_21_3/ab[2][2] ),
	.B(n229),
	.OUT(n228));
   NOR2 U302 (.A(\mult_21_3/ab[4][2] ),
	.B(n231),
	.OUT(n230));
   NOR2 U303 (.A(\mult_21_3/ab[6][2] ),
	.B(n233),
	.OUT(n232));
   NOR2 U304 (.A(\mult_21_3/ab[7][2] ),
	.B(n235),
	.OUT(n234));
   NOR2 U305 (.A(\mult_21_3/ab[2][1] ),
	.B(n237),
	.OUT(n236));
   NOR2 U306 (.A(\mult_21_3/ab[4][1] ),
	.B(n239),
	.OUT(n238));
   NOR2 U307 (.A(\mult_21_3/ab[6][1] ),
	.B(n241),
	.OUT(n240));
   NOR2 U308 (.A(\mult_21_3/ab[7][1] ),
	.B(n243),
	.OUT(n242));
   NOR2 U309 (.A(\mult_21_3/ab[2][0] ),
	.B(n245),
	.OUT(n244));
   NOR2 U310 (.A(\mult_21_3/ab[4][0] ),
	.B(n247),
	.OUT(n246));
   NOR2 U311 (.A(\mult_21_3/ab[6][0] ),
	.B(n249),
	.OUT(n248));
   NOR2 U312 (.A(\mult_21_3/ab[7][0] ),
	.B(n251),
	.OUT(n250));
   NOR2 U313 (.A(\mult_21_3/ab[3][7] ),
	.B(\mult_21_3/ab[4][6] ),
	.OUT(n252));
   NOR2 U314 (.A(\mult_21_3/ab[4][7] ),
	.B(\mult_21_3/ab[5][6] ),
	.OUT(n253));
   NAND2 U315 (.A(n255),
	.B(n256),
	.OUT(n254));
   NOR2 U316 (.A(\mult_21_3/ab[6][7] ),
	.B(\mult_21_3/ab[7][6] ),
	.OUT(n257));
   NOR2 U317 (.A(\mult_21_3/ab[6][5] ),
	.B(n259),
	.OUT(n258));
   NAND2 U318 (.A(n261),
	.B(n262),
	.OUT(n260));
   NOR2 U319 (.A(\mult_21_3/ab[6][4] ),
	.B(n264),
	.OUT(n263));
   NOR2 U320 (.A(\mult_21_3/ab[7][3] ),
	.B(n266),
	.OUT(n265));
   NOR2 U321 (.A(\mult_21_2/ab[1][7] ),
	.B(\mult_21_2/ab[2][6] ),
	.OUT(n267));
   NAND2 U322 (.A(n269),
	.B(n270),
	.OUT(n268));
   NOR2 U323 (.A(\mult_21_2/ab[4][5] ),
	.B(n272),
	.OUT(n271));
   NAND2 U324 (.A(n274),
	.B(n275),
	.OUT(n273));
   NOR2 U325 (.A(\mult_21_2/ab[4][4] ),
	.B(n277),
	.OUT(n276));
   NAND2 U326 (.A(n279),
	.B(n280),
	.OUT(n278));
   NOR2 U327 (.A(\mult_21_2/ab[4][3] ),
	.B(n282),
	.OUT(n281));
   NOR2 U328 (.A(\mult_21_2/ab[6][3] ),
	.B(n284),
	.OUT(n283));
   NOR2 U329 (.A(\mult_21_2/ab[2][2] ),
	.B(n286),
	.OUT(n285));
   NOR2 U330 (.A(\mult_21_2/ab[4][2] ),
	.B(n288),
	.OUT(n287));
   NOR2 U331 (.A(\mult_21_2/ab[6][2] ),
	.B(n290),
	.OUT(n289));
   NOR2 U332 (.A(\mult_21_2/ab[7][2] ),
	.B(n292),
	.OUT(n291));
   NOR2 U333 (.A(\mult_21_2/ab[2][1] ),
	.B(n294),
	.OUT(n293));
   NOR2 U334 (.A(\mult_21_2/ab[4][1] ),
	.B(n296),
	.OUT(n295));
   NOR2 U335 (.A(\mult_21_2/ab[6][1] ),
	.B(n298),
	.OUT(n297));
   NOR2 U336 (.A(\mult_21_2/ab[7][1] ),
	.B(n300),
	.OUT(n299));
   NOR2 U337 (.A(\mult_21_2/ab[2][0] ),
	.B(n302),
	.OUT(n301));
   NOR2 U338 (.A(\mult_21_2/ab[4][0] ),
	.B(n304),
	.OUT(n303));
   NOR2 U339 (.A(\mult_21_2/ab[6][0] ),
	.B(n306),
	.OUT(n305));
   NOR2 U340 (.A(\mult_21_2/ab[7][0] ),
	.B(n308),
	.OUT(n307));
   NOR2 U341 (.A(\mult_21_2/ab[3][7] ),
	.B(\mult_21_2/ab[4][6] ),
	.OUT(n309));
   NOR2 U342 (.A(\mult_21_2/ab[4][7] ),
	.B(\mult_21_2/ab[5][6] ),
	.OUT(n310));
   NAND2 U343 (.A(n312),
	.B(n313),
	.OUT(n311));
   NOR2 U344 (.A(\mult_21_2/ab[6][7] ),
	.B(\mult_21_2/ab[7][6] ),
	.OUT(n314));
   NOR2 U345 (.A(\mult_21_2/ab[6][5] ),
	.B(n316),
	.OUT(n315));
   NAND2 U346 (.A(n318),
	.B(n319),
	.OUT(n317));
   NOR2 U347 (.A(\mult_21_2/ab[6][4] ),
	.B(n321),
	.OUT(n320));
   NOR2 U348 (.A(\mult_21_2/ab[7][3] ),
	.B(n323),
	.OUT(n322));
   NOR2 U349 (.A(\mult_21/ab[1][7] ),
	.B(\mult_21/ab[2][6] ),
	.OUT(n324));
   NAND2 U350 (.A(n326),
	.B(n327),
	.OUT(n325));
   NOR2 U351 (.A(\mult_21/ab[4][5] ),
	.B(n329),
	.OUT(n328));
   NAND2 U352 (.A(n331),
	.B(n332),
	.OUT(n330));
   NOR2 U353 (.A(\mult_21/ab[4][4] ),
	.B(n334),
	.OUT(n333));
   NAND2 U354 (.A(n336),
	.B(n337),
	.OUT(n335));
   NOR2 U355 (.A(\mult_21/ab[4][3] ),
	.B(n339),
	.OUT(n338));
   NOR2 U356 (.A(\mult_21/ab[6][3] ),
	.B(n341),
	.OUT(n340));
   NOR2 U357 (.A(\mult_21/ab[2][2] ),
	.B(n343),
	.OUT(n342));
   NOR2 U358 (.A(\mult_21/ab[4][2] ),
	.B(n345),
	.OUT(n344));
   NOR2 U359 (.A(\mult_21/ab[6][2] ),
	.B(n347),
	.OUT(n346));
   NOR2 U360 (.A(\mult_21/ab[7][2] ),
	.B(n349),
	.OUT(n348));
   NOR2 U361 (.A(\mult_21/ab[2][1] ),
	.B(n351),
	.OUT(n350));
   NOR2 U362 (.A(\mult_21/ab[4][1] ),
	.B(n353),
	.OUT(n352));
   NOR2 U363 (.A(\mult_21/ab[6][1] ),
	.B(n355),
	.OUT(n354));
   NOR2 U364 (.A(\mult_21/ab[7][1] ),
	.B(n357),
	.OUT(n356));
   NOR2 U365 (.A(\mult_21/ab[2][0] ),
	.B(n359),
	.OUT(n358));
   NOR2 U366 (.A(\mult_21/ab[4][0] ),
	.B(n361),
	.OUT(n360));
   NOR2 U367 (.A(\mult_21/ab[6][0] ),
	.B(n363),
	.OUT(n362));
   NOR2 U368 (.A(\mult_21/ab[7][0] ),
	.B(n365),
	.OUT(n364));
   NOR2 U369 (.A(\mult_21/ab[3][7] ),
	.B(\mult_21/ab[4][6] ),
	.OUT(n366));
   NOR2 U370 (.A(\mult_21/ab[4][7] ),
	.B(\mult_21/ab[5][6] ),
	.OUT(n367));
   NAND2 U371 (.A(n369),
	.B(n370),
	.OUT(n368));
   NOR2 U372 (.A(\mult_21/ab[6][7] ),
	.B(\mult_21/ab[7][6] ),
	.OUT(n371));
   NOR2 U373 (.A(\mult_21/ab[6][5] ),
	.B(n373),
	.OUT(n372));
   NAND2 U374 (.A(n375),
	.B(n376),
	.OUT(n374));
   NOR2 U375 (.A(\mult_21/ab[6][4] ),
	.B(n378),
	.OUT(n377));
   NOR2 U376 (.A(\mult_21/ab[7][3] ),
	.B(n380),
	.OUT(n379));
   NOR2 U377 (.A(\mult_20_3/ab[1][7] ),
	.B(\mult_20_3/ab[2][6] ),
	.OUT(n381));
   NAND2 U378 (.A(n383),
	.B(n384),
	.OUT(n382));
   NOR2 U379 (.A(\mult_20_3/ab[4][5] ),
	.B(n386),
	.OUT(n385));
   NAND2 U380 (.A(n388),
	.B(n389),
	.OUT(n387));
   NOR2 U381 (.A(\mult_20_3/ab[4][4] ),
	.B(n391),
	.OUT(n390));
   NAND2 U382 (.A(n393),
	.B(n394),
	.OUT(n392));
   NOR2 U383 (.A(\mult_20_3/ab[4][3] ),
	.B(n396),
	.OUT(n395));
   NOR2 U384 (.A(\mult_20_3/ab[6][3] ),
	.B(n398),
	.OUT(n397));
   NOR2 U385 (.A(\mult_20_3/ab[2][2] ),
	.B(n400),
	.OUT(n399));
   NOR2 U386 (.A(\mult_20_3/ab[4][2] ),
	.B(n402),
	.OUT(n401));
   NOR2 U387 (.A(\mult_20_3/ab[6][2] ),
	.B(n404),
	.OUT(n403));
   NOR2 U388 (.A(\mult_20_3/ab[7][2] ),
	.B(n406),
	.OUT(n405));
   NOR2 U389 (.A(\mult_20_3/ab[2][1] ),
	.B(n408),
	.OUT(n407));
   NOR2 U390 (.A(\mult_20_3/ab[4][1] ),
	.B(n410),
	.OUT(n409));
   NOR2 U391 (.A(\mult_20_3/ab[6][1] ),
	.B(n412),
	.OUT(n411));
   NOR2 U392 (.A(\mult_20_3/ab[7][1] ),
	.B(n414),
	.OUT(n413));
   NOR2 U393 (.A(\mult_20_3/ab[2][0] ),
	.B(n416),
	.OUT(n415));
   NOR2 U394 (.A(\mult_20_3/ab[4][0] ),
	.B(n418),
	.OUT(n417));
   NOR2 U395 (.A(\mult_20_3/ab[6][0] ),
	.B(n420),
	.OUT(n419));
   NOR2 U396 (.A(\mult_20_3/ab[7][0] ),
	.B(n422),
	.OUT(n421));
   NOR2 U397 (.A(\mult_20_3/ab[3][7] ),
	.B(\mult_20_3/ab[4][6] ),
	.OUT(n423));
   NOR2 U398 (.A(\mult_20_3/ab[4][7] ),
	.B(\mult_20_3/ab[5][6] ),
	.OUT(n424));
   NAND2 U399 (.A(n426),
	.B(n427),
	.OUT(n425));
   NOR2 U400 (.A(\mult_20_3/ab[6][7] ),
	.B(\mult_20_3/ab[7][6] ),
	.OUT(n428));
   NOR2 U401 (.A(\mult_20_3/ab[6][5] ),
	.B(n430),
	.OUT(n429));
   NAND2 U402 (.A(n432),
	.B(n433),
	.OUT(n431));
   NOR2 U403 (.A(\mult_20_3/ab[6][4] ),
	.B(n435),
	.OUT(n434));
   NOR2 U404 (.A(\mult_20_3/ab[7][3] ),
	.B(n437),
	.OUT(n436));
   NOR2 U405 (.A(\mult_20_2/ab[1][7] ),
	.B(\mult_20_2/ab[2][6] ),
	.OUT(n438));
   NAND2 U406 (.A(n440),
	.B(n441),
	.OUT(n439));
   NOR2 U407 (.A(\mult_20_2/ab[4][5] ),
	.B(n443),
	.OUT(n442));
   NAND2 U408 (.A(n445),
	.B(n446),
	.OUT(n444));
   NOR2 U409 (.A(\mult_20_2/ab[4][4] ),
	.B(n448),
	.OUT(n447));
   NAND2 U410 (.A(n450),
	.B(n451),
	.OUT(n449));
   NOR2 U411 (.A(\mult_20_2/ab[4][3] ),
	.B(n453),
	.OUT(n452));
   NOR2 U412 (.A(\mult_20_2/ab[6][3] ),
	.B(n455),
	.OUT(n454));
   NOR2 U413 (.A(\mult_20_2/ab[2][2] ),
	.B(n457),
	.OUT(n456));
   NOR2 U414 (.A(\mult_20_2/ab[4][2] ),
	.B(n459),
	.OUT(n458));
   NOR2 U415 (.A(\mult_20_2/ab[6][2] ),
	.B(n461),
	.OUT(n460));
   NOR2 U416 (.A(\mult_20_2/ab[7][2] ),
	.B(n463),
	.OUT(n462));
   NOR2 U417 (.A(\mult_20_2/ab[2][1] ),
	.B(n465),
	.OUT(n464));
   NOR2 U418 (.A(\mult_20_2/ab[4][1] ),
	.B(n467),
	.OUT(n466));
   NOR2 U419 (.A(\mult_20_2/ab[6][1] ),
	.B(n469),
	.OUT(n468));
   NOR2 U420 (.A(\mult_20_2/ab[7][1] ),
	.B(n471),
	.OUT(n470));
   NOR2 U421 (.A(\mult_20_2/ab[2][0] ),
	.B(n473),
	.OUT(n472));
   NOR2 U422 (.A(\mult_20_2/ab[4][0] ),
	.B(n475),
	.OUT(n474));
   NOR2 U423 (.A(\mult_20_2/ab[6][0] ),
	.B(n477),
	.OUT(n476));
   NOR2 U424 (.A(\mult_20_2/ab[7][0] ),
	.B(n479),
	.OUT(n478));
   NOR2 U425 (.A(\mult_20_2/ab[3][7] ),
	.B(\mult_20_2/ab[4][6] ),
	.OUT(n480));
   NOR2 U426 (.A(\mult_20_2/ab[4][7] ),
	.B(\mult_20_2/ab[5][6] ),
	.OUT(n481));
   NAND2 U427 (.A(n483),
	.B(n484),
	.OUT(n482));
   NOR2 U428 (.A(\mult_20_2/ab[6][7] ),
	.B(\mult_20_2/ab[7][6] ),
	.OUT(n485));
   NOR2 U429 (.A(\mult_20_2/ab[6][5] ),
	.B(n487),
	.OUT(n486));
   NAND2 U430 (.A(n489),
	.B(n490),
	.OUT(n488));
   NOR2 U431 (.A(\mult_20_2/ab[6][4] ),
	.B(n492),
	.OUT(n491));
   NOR2 U432 (.A(\mult_20_2/ab[7][3] ),
	.B(n494),
	.OUT(n493));
   NOR2 U433 (.A(\mult_20/ab[1][7] ),
	.B(\mult_20/ab[2][6] ),
	.OUT(n495));
   NAND2 U434 (.A(n497),
	.B(n498),
	.OUT(n496));
   NOR2 U435 (.A(\mult_20/ab[4][5] ),
	.B(n500),
	.OUT(n499));
   NAND2 U436 (.A(n502),
	.B(n503),
	.OUT(n501));
   NOR2 U437 (.A(\mult_20/ab[4][4] ),
	.B(n505),
	.OUT(n504));
   NAND2 U438 (.A(n507),
	.B(n508),
	.OUT(n506));
   NOR2 U439 (.A(\mult_20/ab[4][3] ),
	.B(n510),
	.OUT(n509));
   NOR2 U440 (.A(\mult_20/ab[6][3] ),
	.B(n512),
	.OUT(n511));
   NOR2 U441 (.A(\mult_20/ab[2][2] ),
	.B(n514),
	.OUT(n513));
   NOR2 U442 (.A(\mult_20/ab[4][2] ),
	.B(n516),
	.OUT(n515));
   NOR2 U443 (.A(\mult_20/ab[6][2] ),
	.B(n518),
	.OUT(n517));
   NOR2 U444 (.A(\mult_20/ab[7][2] ),
	.B(n520),
	.OUT(n519));
   NOR2 U445 (.A(\mult_20/ab[2][1] ),
	.B(n522),
	.OUT(n521));
   NOR2 U446 (.A(\mult_20/ab[4][1] ),
	.B(n524),
	.OUT(n523));
   NOR2 U447 (.A(\mult_20/ab[6][1] ),
	.B(n526),
	.OUT(n525));
   NOR2 U448 (.A(\mult_20/ab[7][1] ),
	.B(n528),
	.OUT(n527));
   NOR2 U449 (.A(\mult_20/ab[2][0] ),
	.B(n530),
	.OUT(n529));
   NOR2 U450 (.A(\mult_20/ab[4][0] ),
	.B(n532),
	.OUT(n531));
   NOR2 U451 (.A(\mult_20/ab[6][0] ),
	.B(n534),
	.OUT(n533));
   NOR2 U452 (.A(\mult_20/ab[7][0] ),
	.B(n536),
	.OUT(n535));
   NOR2 U453 (.A(\mult_20/ab[3][7] ),
	.B(\mult_20/ab[4][6] ),
	.OUT(n537));
   NOR2 U454 (.A(\mult_20/ab[4][7] ),
	.B(\mult_20/ab[5][6] ),
	.OUT(n538));
   NAND2 U455 (.A(n540),
	.B(n541),
	.OUT(n539));
   NOR2 U456 (.A(\mult_20/ab[6][7] ),
	.B(\mult_20/ab[7][6] ),
	.OUT(n542));
   NOR2 U457 (.A(\mult_20/ab[6][5] ),
	.B(n544),
	.OUT(n543));
   NAND2 U458 (.A(n546),
	.B(n547),
	.OUT(n545));
   NOR2 U459 (.A(\mult_20/ab[6][4] ),
	.B(n549),
	.OUT(n548));
   NOR2 U460 (.A(\mult_20/ab[7][3] ),
	.B(n551),
	.OUT(n550));
   NOR2 U461 (.A(\mult_19_3/ab[1][7] ),
	.B(\mult_19_3/ab[2][6] ),
	.OUT(n552));
   NAND2 U462 (.A(n554),
	.B(n555),
	.OUT(n553));
   NOR2 U463 (.A(\mult_19_3/ab[4][5] ),
	.B(n557),
	.OUT(n556));
   NAND2 U464 (.A(n559),
	.B(n560),
	.OUT(n558));
   NOR2 U465 (.A(\mult_19_3/ab[4][4] ),
	.B(n562),
	.OUT(n561));
   NAND2 U466 (.A(n564),
	.B(n565),
	.OUT(n563));
   NOR2 U467 (.A(\mult_19_3/ab[4][3] ),
	.B(n567),
	.OUT(n566));
   NOR2 U468 (.A(\mult_19_3/ab[6][3] ),
	.B(n569),
	.OUT(n568));
   NOR2 U469 (.A(\mult_19_3/ab[2][2] ),
	.B(n571),
	.OUT(n570));
   NOR2 U470 (.A(\mult_19_3/ab[4][2] ),
	.B(n573),
	.OUT(n572));
   NOR2 U471 (.A(\mult_19_3/ab[6][2] ),
	.B(n575),
	.OUT(n574));
   NOR2 U472 (.A(\mult_19_3/ab[7][2] ),
	.B(n577),
	.OUT(n576));
   NOR2 U473 (.A(\mult_19_3/ab[2][1] ),
	.B(n579),
	.OUT(n578));
   NOR2 U474 (.A(\mult_19_3/ab[4][1] ),
	.B(n581),
	.OUT(n580));
   NOR2 U475 (.A(\mult_19_3/ab[6][1] ),
	.B(n583),
	.OUT(n582));
   NOR2 U476 (.A(\mult_19_3/ab[7][1] ),
	.B(n585),
	.OUT(n584));
   NOR2 U477 (.A(\mult_19_3/ab[2][0] ),
	.B(n587),
	.OUT(n586));
   NOR2 U478 (.A(\mult_19_3/ab[4][0] ),
	.B(n589),
	.OUT(n588));
   NOR2 U479 (.A(\mult_19_3/ab[6][0] ),
	.B(n591),
	.OUT(n590));
   NOR2 U480 (.A(\mult_19_3/ab[7][0] ),
	.B(n593),
	.OUT(n592));
   NOR2 U481 (.A(\mult_19_3/ab[3][7] ),
	.B(\mult_19_3/ab[4][6] ),
	.OUT(n594));
   NOR2 U482 (.A(\mult_19_3/ab[4][7] ),
	.B(\mult_19_3/ab[5][6] ),
	.OUT(n595));
   NAND2 U483 (.A(n597),
	.B(n598),
	.OUT(n596));
   NOR2 U484 (.A(\mult_19_3/ab[6][7] ),
	.B(\mult_19_3/ab[7][6] ),
	.OUT(n599));
   NOR2 U485 (.A(\mult_19_3/ab[6][5] ),
	.B(n601),
	.OUT(n600));
   NAND2 U486 (.A(n603),
	.B(n604),
	.OUT(n602));
   NOR2 U487 (.A(\mult_19_3/ab[6][4] ),
	.B(n606),
	.OUT(n605));
   NOR2 U488 (.A(\mult_19_3/ab[7][3] ),
	.B(n608),
	.OUT(n607));
   NOR2 U489 (.A(\mult_19_2/ab[1][7] ),
	.B(\mult_19_2/ab[2][6] ),
	.OUT(n609));
   NAND2 U490 (.A(n611),
	.B(n612),
	.OUT(n610));
   NOR2 U491 (.A(\mult_19_2/ab[4][5] ),
	.B(n614),
	.OUT(n613));
   NAND2 U492 (.A(n616),
	.B(n617),
	.OUT(n615));
   NOR2 U493 (.A(\mult_19_2/ab[4][4] ),
	.B(n619),
	.OUT(n618));
   NAND2 U494 (.A(n621),
	.B(n622),
	.OUT(n620));
   NOR2 U495 (.A(\mult_19_2/ab[4][3] ),
	.B(n624),
	.OUT(n623));
   NOR2 U496 (.A(\mult_19_2/ab[6][3] ),
	.B(n626),
	.OUT(n625));
   NOR2 U497 (.A(\mult_19_2/ab[2][2] ),
	.B(n628),
	.OUT(n627));
   NOR2 U498 (.A(\mult_19_2/ab[4][2] ),
	.B(n630),
	.OUT(n629));
   NOR2 U499 (.A(\mult_19_2/ab[6][2] ),
	.B(n632),
	.OUT(n631));
   NOR2 U500 (.A(\mult_19_2/ab[7][2] ),
	.B(n634),
	.OUT(n633));
   NOR2 U501 (.A(\mult_19_2/ab[2][1] ),
	.B(n636),
	.OUT(n635));
   NOR2 U502 (.A(\mult_19_2/ab[4][1] ),
	.B(n638),
	.OUT(n637));
   NOR2 U503 (.A(\mult_19_2/ab[6][1] ),
	.B(n640),
	.OUT(n639));
   NOR2 U504 (.A(\mult_19_2/ab[7][1] ),
	.B(n642),
	.OUT(n641));
   NOR2 U505 (.A(\mult_19_2/ab[2][0] ),
	.B(n644),
	.OUT(n643));
   NOR2 U506 (.A(\mult_19_2/ab[4][0] ),
	.B(n646),
	.OUT(n645));
   NOR2 U507 (.A(\mult_19_2/ab[6][0] ),
	.B(n648),
	.OUT(n647));
   NOR2 U508 (.A(\mult_19_2/ab[7][0] ),
	.B(n650),
	.OUT(n649));
   NOR2 U509 (.A(\mult_19_2/ab[3][7] ),
	.B(\mult_19_2/ab[4][6] ),
	.OUT(n651));
   NOR2 U510 (.A(\mult_19_2/ab[4][7] ),
	.B(\mult_19_2/ab[5][6] ),
	.OUT(n652));
   NAND2 U511 (.A(n654),
	.B(n655),
	.OUT(n653));
   NOR2 U512 (.A(\mult_19_2/ab[6][7] ),
	.B(\mult_19_2/ab[7][6] ),
	.OUT(n656));
   NOR2 U513 (.A(\mult_19_2/ab[6][5] ),
	.B(n658),
	.OUT(n657));
   NAND2 U514 (.A(n660),
	.B(n661),
	.OUT(n659));
   NOR2 U515 (.A(\mult_19_2/ab[6][4] ),
	.B(n663),
	.OUT(n662));
   NOR2 U516 (.A(\mult_19_2/ab[7][3] ),
	.B(n665),
	.OUT(n664));
   NOR2 U517 (.A(\mult_19/ab[1][7] ),
	.B(\mult_19/ab[2][6] ),
	.OUT(n666));
   NAND2 U518 (.A(n668),
	.B(n669),
	.OUT(n667));
   NOR2 U519 (.A(\mult_19/ab[4][5] ),
	.B(n671),
	.OUT(n670));
   NAND2 U520 (.A(n673),
	.B(n674),
	.OUT(n672));
   NOR2 U521 (.A(\mult_19/ab[4][4] ),
	.B(n676),
	.OUT(n675));
   NAND2 U522 (.A(n678),
	.B(n679),
	.OUT(n677));
   NOR2 U523 (.A(\mult_19/ab[4][3] ),
	.B(n681),
	.OUT(n680));
   NOR2 U524 (.A(\mult_19/ab[6][3] ),
	.B(n683),
	.OUT(n682));
   NOR2 U525 (.A(\mult_19/ab[2][2] ),
	.B(n685),
	.OUT(n684));
   NOR2 U526 (.A(\mult_19/ab[4][2] ),
	.B(n687),
	.OUT(n686));
   NOR2 U527 (.A(\mult_19/ab[6][2] ),
	.B(n689),
	.OUT(n688));
   NOR2 U528 (.A(\mult_19/ab[7][2] ),
	.B(n691),
	.OUT(n690));
   NOR2 U529 (.A(\mult_19/ab[2][1] ),
	.B(n693),
	.OUT(n692));
   NOR2 U530 (.A(\mult_19/ab[4][1] ),
	.B(n695),
	.OUT(n694));
   NOR2 U531 (.A(\mult_19/ab[6][1] ),
	.B(n697),
	.OUT(n696));
   NOR2 U532 (.A(\mult_19/ab[7][1] ),
	.B(n699),
	.OUT(n698));
   NOR2 U533 (.A(\mult_19/ab[2][0] ),
	.B(n701),
	.OUT(n700));
   NOR2 U534 (.A(\mult_19/ab[4][0] ),
	.B(n703),
	.OUT(n702));
   NOR2 U535 (.A(\mult_19/ab[6][0] ),
	.B(n705),
	.OUT(n704));
   NOR2 U536 (.A(\mult_19/ab[7][0] ),
	.B(n707),
	.OUT(n706));
   NOR2 U537 (.A(\mult_19/ab[3][7] ),
	.B(\mult_19/ab[4][6] ),
	.OUT(n708));
   NOR2 U538 (.A(\mult_19/ab[4][7] ),
	.B(\mult_19/ab[5][6] ),
	.OUT(n709));
   NAND2 U539 (.A(n711),
	.B(n712),
	.OUT(n710));
   NOR2 U540 (.A(\mult_19/ab[6][7] ),
	.B(\mult_19/ab[7][6] ),
	.OUT(n713));
   NOR2 U541 (.A(\mult_19/ab[6][5] ),
	.B(n715),
	.OUT(n714));
   NAND2 U542 (.A(n717),
	.B(n718),
	.OUT(n716));
   NOR2 U543 (.A(\mult_19/ab[6][4] ),
	.B(n720),
	.OUT(n719));
   NOR2 U544 (.A(\mult_19/ab[7][3] ),
	.B(n722),
	.OUT(n721));
   NOR2 U545 (.A(N20),
	.B(N4),
	.OUT(n723));
   NOR2 U546 (.A(N21),
	.B(N5),
	.OUT(n724));
   NOR2 U547 (.A(N22),
	.B(N6),
	.OUT(n725));
   NOR2 U548 (.A(N23),
	.B(N7),
	.OUT(n726));
   NOR2 U549 (.A(N24),
	.B(N8),
	.OUT(n727));
   NOR2 U550 (.A(N25),
	.B(N9),
	.OUT(n728));
   NOR2 U551 (.A(N26),
	.B(N10),
	.OUT(n729));
   NOR2 U552 (.A(N27),
	.B(N11),
	.OUT(n730));
   NOR2 U553 (.A(N28),
	.B(N12),
	.OUT(n731));
   NOR2 U554 (.A(N29),
	.B(N13),
	.OUT(n732));
   NOR2 U555 (.A(N30),
	.B(N14),
	.OUT(n733));
   NOR2 U556 (.A(N31),
	.B(N15),
	.OUT(n734));
   NOR2 U557 (.A(n736),
	.B(n737),
	.OUT(n735));
   NAND2 U558 (.A(n739),
	.B(n740),
	.OUT(n738));
   NOR2 U559 (.A(N53),
	.B(n742),
	.OUT(n741));
   NAND2 U560 (.A(n744),
	.B(n745),
	.OUT(n743));
   NOR2 U561 (.A(N56),
	.B(n747),
	.OUT(n746));
   NOR2 U562 (.A(N57),
	.B(n749),
	.OUT(n748));
   NAND2 U563 (.A(n751),
	.B(n752),
	.OUT(n750));
   NOR2 U564 (.A(N59),
	.B(n754),
	.OUT(n753));
   NAND2 U565 (.A(n756),
	.B(n757),
	.OUT(n755));
   NOR2 U566 (.A(N61),
	.B(n759),
	.OUT(n758));
   NAND2 U567 (.A(n761),
	.B(n762),
	.OUT(n760));
   NOR2 U568 (.A(N63),
	.B(n764),
	.OUT(n763));
   NOR2 U569 (.A(N180),
	.B(N164),
	.OUT(n765));
   NOR2 U570 (.A(N181),
	.B(N165),
	.OUT(n766));
   NOR2 U571 (.A(N182),
	.B(N166),
	.OUT(n767));
   NOR2 U572 (.A(N183),
	.B(N167),
	.OUT(n768));
   NOR2 U573 (.A(N184),
	.B(N168),
	.OUT(n769));
   NOR2 U574 (.A(N185),
	.B(N169),
	.OUT(n770));
   NOR2 U575 (.A(N186),
	.B(N170),
	.OUT(n771));
   NOR2 U576 (.A(N187),
	.B(N171),
	.OUT(n772));
   NOR2 U577 (.A(N188),
	.B(N172),
	.OUT(n773));
   NOR2 U578 (.A(N189),
	.B(N173),
	.OUT(n774));
   NOR2 U579 (.A(N190),
	.B(N174),
	.OUT(n775));
   NOR2 U580 (.A(N191),
	.B(N175),
	.OUT(n776));
   NOR2 U581 (.A(n778),
	.B(n779),
	.OUT(n777));
   NAND2 U582 (.A(n781),
	.B(n782),
	.OUT(n780));
   NOR2 U583 (.A(N213),
	.B(n784),
	.OUT(n783));
   NAND2 U584 (.A(n786),
	.B(n787),
	.OUT(n785));
   NOR2 U585 (.A(N216),
	.B(n789),
	.OUT(n788));
   NOR2 U586 (.A(N217),
	.B(n791),
	.OUT(n790));
   NAND2 U587 (.A(n793),
	.B(n794),
	.OUT(n792));
   NOR2 U588 (.A(N219),
	.B(n796),
	.OUT(n795));
   NAND2 U589 (.A(n798),
	.B(n799),
	.OUT(n797));
   NOR2 U590 (.A(N221),
	.B(n801),
	.OUT(n800));
   NAND2 U591 (.A(n803),
	.B(n804),
	.OUT(n802));
   NOR2 U592 (.A(N223),
	.B(n806),
	.OUT(n805));
   NOR2 U593 (.A(N100),
	.B(N84),
	.OUT(n807));
   NOR2 U594 (.A(N101),
	.B(N85),
	.OUT(n808));
   NOR2 U595 (.A(N102),
	.B(N86),
	.OUT(n809));
   NOR2 U596 (.A(N103),
	.B(N87),
	.OUT(n810));
   NOR2 U597 (.A(N104),
	.B(N88),
	.OUT(n811));
   NOR2 U598 (.A(N105),
	.B(N89),
	.OUT(n812));
   NOR2 U599 (.A(N106),
	.B(N90),
	.OUT(n813));
   NOR2 U600 (.A(N107),
	.B(N91),
	.OUT(n814));
   NOR2 U601 (.A(N108),
	.B(N92),
	.OUT(n815));
   NOR2 U602 (.A(N109),
	.B(N93),
	.OUT(n816));
   NOR2 U603 (.A(N110),
	.B(N94),
	.OUT(n817));
   NOR2 U604 (.A(N111),
	.B(N95),
	.OUT(n818));
   NOR2 U605 (.A(n820),
	.B(n821),
	.OUT(n819));
   NAND2 U606 (.A(n823),
	.B(n824),
	.OUT(n822));
   NOR2 U607 (.A(N133),
	.B(n826),
	.OUT(n825));
   NAND2 U608 (.A(n828),
	.B(n829),
	.OUT(n827));
   NOR2 U609 (.A(N136),
	.B(n831),
	.OUT(n830));
   NOR2 U610 (.A(N137),
	.B(n833),
	.OUT(n832));
   NAND2 U611 (.A(n835),
	.B(n836),
	.OUT(n834));
   NOR2 U612 (.A(N139),
	.B(n838),
	.OUT(n837));
   NAND2 U613 (.A(n840),
	.B(n841),
	.OUT(n839));
   NOR2 U614 (.A(N141),
	.B(n843),
	.OUT(n842));
   NAND2 U615 (.A(n845),
	.B(n846),
	.OUT(n844));
   NOR2 U616 (.A(N143),
	.B(n848),
	.OUT(n847));
   XOR2 U617 (.A(\mult_21_3/ab[1][7] ),
	.B(n850),
	.OUT(n849));
   XOR2 U618 (.A(\mult_21_3/ab[1][6] ),
	.B(\mult_21_3/ab[0][7] ),
	.OUT(n851));
   XOR2 U619 (.A(\mult_21_3/ab[1][5] ),
	.B(\mult_21_3/ab[0][6] ),
	.OUT(n852));
   XOR2 U620 (.A(n851),
	.B(n854),
	.OUT(n853));
   XOR2 U621 (.A(n856),
	.B(n857),
	.OUT(n855));
   XOR2 U622 (.A(\mult_21_3/ab[1][4] ),
	.B(\mult_21_3/ab[0][5] ),
	.OUT(n858));
   XOR2 U623 (.A(n852),
	.B(n860),
	.OUT(n859));
   XOR2 U624 (.A(\mult_21_3/ab[1][3] ),
	.B(\mult_21_3/ab[0][4] ),
	.OUT(n861));
   XOR2 U625 (.A(n858),
	.B(n863),
	.OUT(n862));
   XOR2 U626 (.A(n865),
	.B(n866),
	.OUT(n864));
   XOR2 U627 (.A(n868),
	.B(n869),
	.OUT(n867));
   XOR2 U628 (.A(n871),
	.B(n872),
	.OUT(n870));
   XOR2 U629 (.A(n874),
	.B(n875),
	.OUT(n873));
   XOR2 U630 (.A(n876),
	.B(n877),
	.OUT(n205));
   XOR2 U631 (.A(\mult_21_3/ab[1][2] ),
	.B(\mult_21_3/ab[0][3] ),
	.OUT(n878));
   XOR2 U632 (.A(n861),
	.B(n880),
	.OUT(n879));
   XOR2 U633 (.A(n882),
	.B(n883),
	.OUT(n881));
   XOR2 U634 (.A(n885),
	.B(n886),
	.OUT(n884));
   XOR2 U635 (.A(\mult_21_3/ab[1][1] ),
	.B(\mult_21_3/ab[0][2] ),
	.OUT(n887));
   XOR2 U636 (.A(n878),
	.B(n889),
	.OUT(n888));
   XOR2 U637 (.A(n891),
	.B(n892),
	.OUT(n890));
   XOR2 U638 (.A(n894),
	.B(n895),
	.OUT(n893));
   XOR2 U639 (.A(n897),
	.B(n898),
	.OUT(n896));
   XOR2 U640 (.A(n899),
	.B(n900),
	.OUT(n201));
   XOR2 U641 (.A(n204),
	.B(n205),
	.OUT(\mult_21_3/A1[8] ));
   XOR2 U642 (.A(n901),
	.B(n902),
	.OUT(\mult_21_3/A1[5] ));
   XOR2 U643 (.A(n890),
	.B(n903),
	.OUT(\mult_21_3/A1[3] ));
   XOR2 U644 (.A(n888),
	.B(n905),
	.OUT(n904));
   XOR2 U645 (.A(n195),
	.B(n194),
	.OUT(\mult_21_3/A1[12] ));
   XOR2 U646 (.A(n200),
	.B(n201),
	.OUT(\mult_21_3/A1[10] ));
   XOR2 U647 (.A(\mult_21_2/ab[1][7] ),
	.B(n907),
	.OUT(n906));
   XOR2 U648 (.A(\mult_21_2/ab[1][6] ),
	.B(\mult_21_2/ab[0][7] ),
	.OUT(n908));
   XOR2 U649 (.A(\mult_21_2/ab[1][5] ),
	.B(\mult_21_2/ab[0][6] ),
	.OUT(n909));
   XOR2 U650 (.A(n908),
	.B(n911),
	.OUT(n910));
   XOR2 U651 (.A(n913),
	.B(n914),
	.OUT(n912));
   XOR2 U652 (.A(\mult_21_2/ab[1][4] ),
	.B(\mult_21_2/ab[0][5] ),
	.OUT(n915));
   XOR2 U653 (.A(n909),
	.B(n917),
	.OUT(n916));
   XOR2 U654 (.A(\mult_21_2/ab[1][3] ),
	.B(\mult_21_2/ab[0][4] ),
	.OUT(n918));
   XOR2 U655 (.A(n915),
	.B(n920),
	.OUT(n919));
   XOR2 U656 (.A(n922),
	.B(n923),
	.OUT(n921));
   XOR2 U657 (.A(n925),
	.B(n926),
	.OUT(n924));
   XOR2 U658 (.A(n928),
	.B(n929),
	.OUT(n927));
   XOR2 U659 (.A(n931),
	.B(n932),
	.OUT(n930));
   XOR2 U660 (.A(n933),
	.B(n934),
	.OUT(n189));
   XOR2 U661 (.A(\mult_21_2/ab[1][2] ),
	.B(\mult_21_2/ab[0][3] ),
	.OUT(n935));
   XOR2 U662 (.A(n918),
	.B(n937),
	.OUT(n936));
   XOR2 U663 (.A(n939),
	.B(n940),
	.OUT(n938));
   XOR2 U664 (.A(n942),
	.B(n943),
	.OUT(n941));
   XOR2 U665 (.A(\mult_21_2/ab[1][1] ),
	.B(\mult_21_2/ab[0][2] ),
	.OUT(n944));
   XOR2 U666 (.A(n935),
	.B(n946),
	.OUT(n945));
   XOR2 U667 (.A(n948),
	.B(n949),
	.OUT(n947));
   XOR2 U668 (.A(n951),
	.B(n952),
	.OUT(n950));
   XOR2 U669 (.A(n954),
	.B(n955),
	.OUT(n953));
   XOR2 U670 (.A(n956),
	.B(n957),
	.OUT(n185));
   XOR2 U671 (.A(n188),
	.B(n189),
	.OUT(\mult_21_2/A1[8] ));
   XOR2 U672 (.A(n958),
	.B(n959),
	.OUT(\mult_21_2/A1[5] ));
   XOR2 U673 (.A(n947),
	.B(n960),
	.OUT(\mult_21_2/A1[3] ));
   XOR2 U674 (.A(n945),
	.B(n962),
	.OUT(n961));
   XOR2 U675 (.A(n179),
	.B(n178),
	.OUT(\mult_21_2/A1[12] ));
   XOR2 U676 (.A(n184),
	.B(n185),
	.OUT(\mult_21_2/A1[10] ));
   XOR2 U677 (.A(\mult_21/ab[1][7] ),
	.B(n964),
	.OUT(n963));
   XOR2 U678 (.A(\mult_21/ab[1][6] ),
	.B(\mult_21/ab[0][7] ),
	.OUT(n965));
   XOR2 U679 (.A(\mult_21/ab[1][5] ),
	.B(\mult_21/ab[0][6] ),
	.OUT(n966));
   XOR2 U680 (.A(n965),
	.B(n968),
	.OUT(n967));
   XOR2 U681 (.A(n970),
	.B(n971),
	.OUT(n969));
   XOR2 U682 (.A(\mult_21/ab[1][4] ),
	.B(\mult_21/ab[0][5] ),
	.OUT(n972));
   XOR2 U683 (.A(n966),
	.B(n974),
	.OUT(n973));
   XOR2 U684 (.A(\mult_21/ab[1][3] ),
	.B(\mult_21/ab[0][4] ),
	.OUT(n975));
   XOR2 U685 (.A(n972),
	.B(n977),
	.OUT(n976));
   XOR2 U686 (.A(n979),
	.B(n980),
	.OUT(n978));
   XOR2 U687 (.A(n982),
	.B(n983),
	.OUT(n981));
   XOR2 U688 (.A(n985),
	.B(n986),
	.OUT(n984));
   XOR2 U689 (.A(n988),
	.B(n989),
	.OUT(n987));
   XOR2 U690 (.A(n990),
	.B(n991),
	.OUT(n173));
   XOR2 U691 (.A(\mult_21/ab[1][2] ),
	.B(\mult_21/ab[0][3] ),
	.OUT(n992));
   XOR2 U692 (.A(n975),
	.B(n994),
	.OUT(n993));
   XOR2 U693 (.A(n996),
	.B(n997),
	.OUT(n995));
   XOR2 U694 (.A(n999),
	.B(n1000),
	.OUT(n998));
   XOR2 U695 (.A(\mult_21/ab[1][1] ),
	.B(\mult_21/ab[0][2] ),
	.OUT(n1001));
   XOR2 U696 (.A(n992),
	.B(n1003),
	.OUT(n1002));
   XOR2 U697 (.A(n1005),
	.B(n1006),
	.OUT(n1004));
   XOR2 U698 (.A(n1008),
	.B(n1009),
	.OUT(n1007));
   XOR2 U699 (.A(n1011),
	.B(n1012),
	.OUT(n1010));
   XOR2 U700 (.A(n1013),
	.B(n1014),
	.OUT(n169));
   XOR2 U701 (.A(n172),
	.B(n173),
	.OUT(\mult_21/A1[8] ));
   XOR2 U702 (.A(n1015),
	.B(n1016),
	.OUT(\mult_21/A1[5] ));
   XOR2 U703 (.A(n1004),
	.B(n1017),
	.OUT(\mult_21/A1[3] ));
   XOR2 U704 (.A(n1002),
	.B(n1019),
	.OUT(n1018));
   XOR2 U705 (.A(n163),
	.B(n162),
	.OUT(\mult_21/A1[12] ));
   XOR2 U706 (.A(n168),
	.B(n169),
	.OUT(\mult_21/A1[10] ));
   XOR2 U707 (.A(\mult_20_3/ab[1][7] ),
	.B(n1021),
	.OUT(n1020));
   XOR2 U708 (.A(\mult_20_3/ab[1][6] ),
	.B(\mult_20_3/ab[0][7] ),
	.OUT(n1022));
   XOR2 U709 (.A(\mult_20_3/ab[1][5] ),
	.B(\mult_20_3/ab[0][6] ),
	.OUT(n1023));
   XOR2 U710 (.A(n1022),
	.B(n1025),
	.OUT(n1024));
   XOR2 U711 (.A(n1027),
	.B(n1028),
	.OUT(n1026));
   XOR2 U712 (.A(\mult_20_3/ab[1][4] ),
	.B(\mult_20_3/ab[0][5] ),
	.OUT(n1029));
   XOR2 U713 (.A(n1023),
	.B(n1031),
	.OUT(n1030));
   XOR2 U714 (.A(\mult_20_3/ab[1][3] ),
	.B(\mult_20_3/ab[0][4] ),
	.OUT(n1032));
   XOR2 U715 (.A(n1029),
	.B(n1034),
	.OUT(n1033));
   XOR2 U716 (.A(n1036),
	.B(n1037),
	.OUT(n1035));
   XOR2 U717 (.A(n1039),
	.B(n1040),
	.OUT(n1038));
   XOR2 U718 (.A(n1042),
	.B(n1043),
	.OUT(n1041));
   XOR2 U719 (.A(n1045),
	.B(n1046),
	.OUT(n1044));
   XOR2 U720 (.A(n1047),
	.B(n1048),
	.OUT(n157));
   XOR2 U721 (.A(\mult_20_3/ab[1][2] ),
	.B(\mult_20_3/ab[0][3] ),
	.OUT(n1049));
   XOR2 U722 (.A(n1032),
	.B(n1051),
	.OUT(n1050));
   XOR2 U723 (.A(n1053),
	.B(n1054),
	.OUT(n1052));
   XOR2 U724 (.A(n1056),
	.B(n1057),
	.OUT(n1055));
   XOR2 U725 (.A(\mult_20_3/ab[1][1] ),
	.B(\mult_20_3/ab[0][2] ),
	.OUT(n1058));
   XOR2 U726 (.A(n1049),
	.B(n1060),
	.OUT(n1059));
   XOR2 U727 (.A(n1062),
	.B(n1063),
	.OUT(n1061));
   XOR2 U728 (.A(n1065),
	.B(n1066),
	.OUT(n1064));
   XOR2 U729 (.A(n1068),
	.B(n1069),
	.OUT(n1067));
   XOR2 U730 (.A(n1070),
	.B(n1071),
	.OUT(n153));
   XOR2 U731 (.A(n156),
	.B(n157),
	.OUT(\mult_20_3/A1[8] ));
   XOR2 U732 (.A(n1072),
	.B(n1073),
	.OUT(\mult_20_3/A1[5] ));
   XOR2 U733 (.A(n1061),
	.B(n1074),
	.OUT(\mult_20_3/A1[3] ));
   XOR2 U734 (.A(n1059),
	.B(n1076),
	.OUT(n1075));
   XOR2 U735 (.A(n147),
	.B(n146),
	.OUT(\mult_20_3/A1[12] ));
   XOR2 U736 (.A(n152),
	.B(n153),
	.OUT(\mult_20_3/A1[10] ));
   XOR2 U737 (.A(\mult_20_2/ab[1][7] ),
	.B(n1078),
	.OUT(n1077));
   XOR2 U738 (.A(\mult_20_2/ab[1][6] ),
	.B(\mult_20_2/ab[0][7] ),
	.OUT(n1079));
   XOR2 U739 (.A(\mult_20_2/ab[1][5] ),
	.B(\mult_20_2/ab[0][6] ),
	.OUT(n1080));
   XOR2 U740 (.A(n1079),
	.B(n1082),
	.OUT(n1081));
   XOR2 U741 (.A(n1084),
	.B(n1085),
	.OUT(n1083));
   XOR2 U742 (.A(\mult_20_2/ab[1][4] ),
	.B(\mult_20_2/ab[0][5] ),
	.OUT(n1086));
   XOR2 U743 (.A(n1080),
	.B(n1088),
	.OUT(n1087));
   XOR2 U744 (.A(\mult_20_2/ab[1][3] ),
	.B(\mult_20_2/ab[0][4] ),
	.OUT(n1089));
   XOR2 U745 (.A(n1086),
	.B(n1091),
	.OUT(n1090));
   XOR2 U746 (.A(n1093),
	.B(n1094),
	.OUT(n1092));
   XOR2 U747 (.A(n1096),
	.B(n1097),
	.OUT(n1095));
   XOR2 U748 (.A(n1099),
	.B(n1100),
	.OUT(n1098));
   XOR2 U749 (.A(n1102),
	.B(n1103),
	.OUT(n1101));
   XOR2 U750 (.A(n1104),
	.B(n1105),
	.OUT(n141));
   XOR2 U751 (.A(\mult_20_2/ab[1][2] ),
	.B(\mult_20_2/ab[0][3] ),
	.OUT(n1106));
   XOR2 U752 (.A(n1089),
	.B(n1108),
	.OUT(n1107));
   XOR2 U753 (.A(n1110),
	.B(n1111),
	.OUT(n1109));
   XOR2 U754 (.A(n1113),
	.B(n1114),
	.OUT(n1112));
   XOR2 U755 (.A(\mult_20_2/ab[1][1] ),
	.B(\mult_20_2/ab[0][2] ),
	.OUT(n1115));
   XOR2 U756 (.A(n1106),
	.B(n1117),
	.OUT(n1116));
   XOR2 U757 (.A(n1119),
	.B(n1120),
	.OUT(n1118));
   XOR2 U758 (.A(n1122),
	.B(n1123),
	.OUT(n1121));
   XOR2 U759 (.A(n1125),
	.B(n1126),
	.OUT(n1124));
   XOR2 U760 (.A(n1127),
	.B(n1128),
	.OUT(n137));
   XOR2 U761 (.A(n140),
	.B(n141),
	.OUT(\mult_20_2/A1[8] ));
   XOR2 U762 (.A(n1129),
	.B(n1130),
	.OUT(\mult_20_2/A1[5] ));
   XOR2 U763 (.A(n1118),
	.B(n1131),
	.OUT(\mult_20_2/A1[3] ));
   XOR2 U764 (.A(n1116),
	.B(n1133),
	.OUT(n1132));
   XOR2 U765 (.A(n131),
	.B(n130),
	.OUT(\mult_20_2/A1[12] ));
   XOR2 U766 (.A(n136),
	.B(n137),
	.OUT(\mult_20_2/A1[10] ));
   XOR2 U767 (.A(\mult_20/ab[1][7] ),
	.B(n1135),
	.OUT(n1134));
   XOR2 U768 (.A(\mult_20/ab[1][6] ),
	.B(\mult_20/ab[0][7] ),
	.OUT(n1136));
   XOR2 U769 (.A(\mult_20/ab[1][5] ),
	.B(\mult_20/ab[0][6] ),
	.OUT(n1137));
   XOR2 U770 (.A(n1136),
	.B(n1139),
	.OUT(n1138));
   XOR2 U771 (.A(n1141),
	.B(n1142),
	.OUT(n1140));
   XOR2 U772 (.A(\mult_20/ab[1][4] ),
	.B(\mult_20/ab[0][5] ),
	.OUT(n1143));
   XOR2 U773 (.A(n1137),
	.B(n1145),
	.OUT(n1144));
   XOR2 U774 (.A(\mult_20/ab[1][3] ),
	.B(\mult_20/ab[0][4] ),
	.OUT(n1146));
   XOR2 U775 (.A(n1143),
	.B(n1148),
	.OUT(n1147));
   XOR2 U776 (.A(n1150),
	.B(n1151),
	.OUT(n1149));
   XOR2 U777 (.A(n1153),
	.B(n1154),
	.OUT(n1152));
   XOR2 U778 (.A(n1156),
	.B(n1157),
	.OUT(n1155));
   XOR2 U779 (.A(n1159),
	.B(n1160),
	.OUT(n1158));
   XOR2 U780 (.A(n1161),
	.B(n1162),
	.OUT(n125));
   XOR2 U781 (.A(\mult_20/ab[1][2] ),
	.B(\mult_20/ab[0][3] ),
	.OUT(n1163));
   XOR2 U782 (.A(n1146),
	.B(n1165),
	.OUT(n1164));
   XOR2 U783 (.A(n1167),
	.B(n1168),
	.OUT(n1166));
   XOR2 U784 (.A(n1170),
	.B(n1171),
	.OUT(n1169));
   XOR2 U785 (.A(\mult_20/ab[1][1] ),
	.B(\mult_20/ab[0][2] ),
	.OUT(n1172));
   XOR2 U786 (.A(n1163),
	.B(n1174),
	.OUT(n1173));
   XOR2 U787 (.A(n1176),
	.B(n1177),
	.OUT(n1175));
   XOR2 U788 (.A(n1179),
	.B(n1180),
	.OUT(n1178));
   XOR2 U789 (.A(n1182),
	.B(n1183),
	.OUT(n1181));
   XOR2 U790 (.A(n1184),
	.B(n1185),
	.OUT(n121));
   XOR2 U791 (.A(n124),
	.B(n125),
	.OUT(\mult_20/A1[8] ));
   XOR2 U792 (.A(n1186),
	.B(n1187),
	.OUT(\mult_20/A1[5] ));
   XOR2 U793 (.A(n1175),
	.B(n1188),
	.OUT(\mult_20/A1[3] ));
   XOR2 U794 (.A(n1173),
	.B(n1190),
	.OUT(n1189));
   XOR2 U795 (.A(n115),
	.B(n114),
	.OUT(\mult_20/A1[12] ));
   XOR2 U796 (.A(n120),
	.B(n121),
	.OUT(\mult_20/A1[10] ));
   XOR2 U797 (.A(\mult_19_3/ab[1][7] ),
	.B(n1192),
	.OUT(n1191));
   XOR2 U798 (.A(\mult_19_3/ab[1][6] ),
	.B(\mult_19_3/ab[0][7] ),
	.OUT(n1193));
   XOR2 U799 (.A(\mult_19_3/ab[1][5] ),
	.B(\mult_19_3/ab[0][6] ),
	.OUT(n1194));
   XOR2 U800 (.A(n1193),
	.B(n1196),
	.OUT(n1195));
   XOR2 U801 (.A(n1198),
	.B(n1199),
	.OUT(n1197));
   XOR2 U802 (.A(\mult_19_3/ab[1][4] ),
	.B(\mult_19_3/ab[0][5] ),
	.OUT(n1200));
   XOR2 U803 (.A(n1194),
	.B(n1202),
	.OUT(n1201));
   XOR2 U804 (.A(\mult_19_3/ab[1][3] ),
	.B(\mult_19_3/ab[0][4] ),
	.OUT(n1203));
   XOR2 U805 (.A(n1200),
	.B(n1205),
	.OUT(n1204));
   XOR2 U806 (.A(n1207),
	.B(n1208),
	.OUT(n1206));
   XOR2 U807 (.A(n1210),
	.B(n1211),
	.OUT(n1209));
   XOR2 U808 (.A(n1213),
	.B(n1214),
	.OUT(n1212));
   XOR2 U809 (.A(n1216),
	.B(n1217),
	.OUT(n1215));
   XOR2 U810 (.A(n1218),
	.B(n1219),
	.OUT(n109));
   XOR2 U811 (.A(\mult_19_3/ab[1][2] ),
	.B(\mult_19_3/ab[0][3] ),
	.OUT(n1220));
   XOR2 U812 (.A(n1203),
	.B(n1222),
	.OUT(n1221));
   XOR2 U813 (.A(n1224),
	.B(n1225),
	.OUT(n1223));
   XOR2 U814 (.A(n1227),
	.B(n1228),
	.OUT(n1226));
   XOR2 U815 (.A(\mult_19_3/ab[1][1] ),
	.B(\mult_19_3/ab[0][2] ),
	.OUT(n1229));
   XOR2 U816 (.A(n1220),
	.B(n1231),
	.OUT(n1230));
   XOR2 U817 (.A(n1233),
	.B(n1234),
	.OUT(n1232));
   XOR2 U818 (.A(n1236),
	.B(n1237),
	.OUT(n1235));
   XOR2 U819 (.A(n1239),
	.B(n1240),
	.OUT(n1238));
   XOR2 U820 (.A(n1241),
	.B(n1242),
	.OUT(n105));
   XOR2 U821 (.A(n108),
	.B(n109),
	.OUT(\mult_19_3/A1[8] ));
   XOR2 U822 (.A(n1243),
	.B(n1244),
	.OUT(\mult_19_3/A1[5] ));
   XOR2 U823 (.A(n1232),
	.B(n1245),
	.OUT(\mult_19_3/A1[3] ));
   XOR2 U824 (.A(n1230),
	.B(n1247),
	.OUT(n1246));
   XOR2 U825 (.A(n99),
	.B(n98),
	.OUT(\mult_19_3/A1[12] ));
   XOR2 U826 (.A(n104),
	.B(n105),
	.OUT(\mult_19_3/A1[10] ));
   XOR2 U827 (.A(\mult_19_2/ab[1][7] ),
	.B(n1249),
	.OUT(n1248));
   XOR2 U828 (.A(\mult_19_2/ab[1][6] ),
	.B(\mult_19_2/ab[0][7] ),
	.OUT(n1250));
   XOR2 U829 (.A(\mult_19_2/ab[1][5] ),
	.B(\mult_19_2/ab[0][6] ),
	.OUT(n1251));
   XOR2 U830 (.A(n1250),
	.B(n1253),
	.OUT(n1252));
   XOR2 U831 (.A(n1255),
	.B(n1256),
	.OUT(n1254));
   XOR2 U832 (.A(\mult_19_2/ab[1][4] ),
	.B(\mult_19_2/ab[0][5] ),
	.OUT(n1257));
   XOR2 U833 (.A(n1251),
	.B(n1259),
	.OUT(n1258));
   XOR2 U834 (.A(\mult_19_2/ab[1][3] ),
	.B(\mult_19_2/ab[0][4] ),
	.OUT(n1260));
   XOR2 U835 (.A(n1257),
	.B(n1262),
	.OUT(n1261));
   XOR2 U836 (.A(n1264),
	.B(n1265),
	.OUT(n1263));
   XOR2 U837 (.A(n1267),
	.B(n1268),
	.OUT(n1266));
   XOR2 U838 (.A(n1270),
	.B(n1271),
	.OUT(n1269));
   XOR2 U839 (.A(n1273),
	.B(n1274),
	.OUT(n1272));
   XOR2 U840 (.A(n1275),
	.B(n1276),
	.OUT(n93));
   XOR2 U841 (.A(\mult_19_2/ab[1][2] ),
	.B(\mult_19_2/ab[0][3] ),
	.OUT(n1277));
   XOR2 U842 (.A(n1260),
	.B(n1279),
	.OUT(n1278));
   XOR2 U843 (.A(n1281),
	.B(n1282),
	.OUT(n1280));
   XOR2 U844 (.A(n1284),
	.B(n1285),
	.OUT(n1283));
   XOR2 U845 (.A(\mult_19_2/ab[1][1] ),
	.B(\mult_19_2/ab[0][2] ),
	.OUT(n1286));
   XOR2 U846 (.A(n1277),
	.B(n1288),
	.OUT(n1287));
   XOR2 U847 (.A(n1290),
	.B(n1291),
	.OUT(n1289));
   XOR2 U848 (.A(n1293),
	.B(n1294),
	.OUT(n1292));
   XOR2 U849 (.A(n1296),
	.B(n1297),
	.OUT(n1295));
   XOR2 U850 (.A(n1298),
	.B(n1299),
	.OUT(n89));
   XOR2 U851 (.A(n92),
	.B(n93),
	.OUT(\mult_19_2/A1[8] ));
   XOR2 U852 (.A(n1300),
	.B(n1301),
	.OUT(\mult_19_2/A1[5] ));
   XOR2 U853 (.A(n1289),
	.B(n1302),
	.OUT(\mult_19_2/A1[3] ));
   XOR2 U854 (.A(n1287),
	.B(n1304),
	.OUT(n1303));
   XOR2 U855 (.A(n83),
	.B(n82),
	.OUT(\mult_19_2/A1[12] ));
   XOR2 U856 (.A(n88),
	.B(n89),
	.OUT(\mult_19_2/A1[10] ));
   XOR2 U857 (.A(\mult_19/ab[1][7] ),
	.B(n1306),
	.OUT(n1305));
   XOR2 U858 (.A(\mult_19/ab[1][6] ),
	.B(\mult_19/ab[0][7] ),
	.OUT(n1307));
   XOR2 U859 (.A(\mult_19/ab[1][5] ),
	.B(\mult_19/ab[0][6] ),
	.OUT(n1308));
   XOR2 U860 (.A(n1307),
	.B(n1310),
	.OUT(n1309));
   XOR2 U861 (.A(n1312),
	.B(n1313),
	.OUT(n1311));
   XOR2 U862 (.A(\mult_19/ab[1][4] ),
	.B(\mult_19/ab[0][5] ),
	.OUT(n1314));
   XOR2 U863 (.A(n1308),
	.B(n1316),
	.OUT(n1315));
   XOR2 U864 (.A(\mult_19/ab[1][3] ),
	.B(\mult_19/ab[0][4] ),
	.OUT(n1317));
   XOR2 U865 (.A(n1314),
	.B(n1319),
	.OUT(n1318));
   XOR2 U866 (.A(n1321),
	.B(n1322),
	.OUT(n1320));
   XOR2 U867 (.A(n1324),
	.B(n1325),
	.OUT(n1323));
   XOR2 U868 (.A(n1327),
	.B(n1328),
	.OUT(n1326));
   XOR2 U869 (.A(n1330),
	.B(n1331),
	.OUT(n1329));
   XOR2 U870 (.A(n1332),
	.B(n1333),
	.OUT(n77));
   XOR2 U871 (.A(\mult_19/ab[1][2] ),
	.B(\mult_19/ab[0][3] ),
	.OUT(n1334));
   XOR2 U872 (.A(n1317),
	.B(n1336),
	.OUT(n1335));
   XOR2 U873 (.A(n1338),
	.B(n1339),
	.OUT(n1337));
   XOR2 U874 (.A(n1341),
	.B(n1342),
	.OUT(n1340));
   XOR2 U875 (.A(\mult_19/ab[1][1] ),
	.B(\mult_19/ab[0][2] ),
	.OUT(n1343));
   XOR2 U876 (.A(n1334),
	.B(n1345),
	.OUT(n1344));
   XOR2 U877 (.A(n1347),
	.B(n1348),
	.OUT(n1346));
   XOR2 U878 (.A(n1350),
	.B(n1351),
	.OUT(n1349));
   XOR2 U879 (.A(n1353),
	.B(n1354),
	.OUT(n1352));
   XOR2 U880 (.A(n1355),
	.B(n1356),
	.OUT(n73));
   XOR2 U881 (.A(n76),
	.B(n77),
	.OUT(\mult_19/A1[8] ));
   XOR2 U882 (.A(n1357),
	.B(n1358),
	.OUT(\mult_19/A1[5] ));
   XOR2 U883 (.A(n1346),
	.B(n1359),
	.OUT(\mult_19/A1[3] ));
   XOR2 U884 (.A(n1344),
	.B(n1361),
	.OUT(n1360));
   XOR2 U885 (.A(n67),
	.B(n66),
	.OUT(\mult_19/A1[12] ));
   XOR2 U886 (.A(n72),
	.B(n73),
	.OUT(\mult_19/A1[10] ));
   XOR2 U887 (.A(\mult_19_2/ab[1][0] ),
	.B(\mult_19_2/ab[0][1] ),
	.OUT(n1362));
   XOR2 U888 (.A(\mult_19/ab[1][0] ),
	.B(\mult_19/ab[0][1] ),
	.OUT(n1363));
   XOR2 U889 (.A(N17),
	.B(N1),
	.OUT(n1364));
   XOR2 U890 (.A(\mult_19_3/ab[1][0] ),
	.B(\mult_19_3/ab[0][1] ),
	.OUT(n737));
   XOR2 U891 (.A(n1363),
	.B(n1366),
	.OUT(n1365));
   XOR2 U892 (.A(\mult_21_2/ab[1][0] ),
	.B(\mult_21_2/ab[0][1] ),
	.OUT(n1367));
   XOR2 U893 (.A(\mult_21/ab[1][0] ),
	.B(\mult_21/ab[0][1] ),
	.OUT(n1368));
   XOR2 U894 (.A(N177),
	.B(N161),
	.OUT(n1369));
   XOR2 U895 (.A(\mult_21_3/ab[1][0] ),
	.B(\mult_21_3/ab[0][1] ),
	.OUT(n779));
   XOR2 U896 (.A(n1368),
	.B(n1371),
	.OUT(n1370));
   XOR2 U897 (.A(\mult_20_2/ab[1][0] ),
	.B(\mult_20_2/ab[0][1] ),
	.OUT(n1372));
   XOR2 U898 (.A(\mult_20/ab[1][0] ),
	.B(\mult_20/ab[0][1] ),
	.OUT(n1373));
   XOR2 U899 (.A(N97),
	.B(N81),
	.OUT(n1374));
   XOR2 U900 (.A(\mult_20_3/ab[1][0] ),
	.B(\mult_20_3/ab[0][1] ),
	.OUT(n821));
   XOR2 U901 (.A(n1373),
	.B(n1376),
	.OUT(n1375));
   NAND2 U902 (.A(\mult_21_3/ab[0][3] ),
	.B(\mult_21_3/ab[1][2] ),
	.OUT(n1377));
   AOI22 U903 (.A(\mult_21_3/ab[2][2] ),
	.B(n229),
	.C(n1379),
	.D(n861),
	.OUT(n1378));
   NAND2 U904 (.A(\mult_21_3/ab[1][3] ),
	.B(\mult_21_3/ab[0][4] ),
	.OUT(n223));
   INVERTER U905 (.IN(\mult_21_3/ab[3][2] ),
	.OUT(n1380));
   OAI21 U906 (.OUT(n231),
	.C(n1381),
	.B(n1380),
	.A(n1378));
   NAND2 U907 (.A(\mult_21_3/ab[1][4] ),
	.B(\mult_21_3/ab[0][5] ),
	.OUT(n218));
   INVERTER U908 (.IN(\mult_21_3/ab[3][3] ),
	.OUT(n1382));
   AOI22 U909 (.A(n1384),
	.B(\mult_21_3/ab[2][3] ),
	.C(n221),
	.D(n858),
	.OUT(n1383));
   AOI22 U910 (.A(n231),
	.B(\mult_21_3/ab[4][2] ),
	.C(n1386),
	.D(n882),
	.OUT(n1385));
   NAND2 U911 (.A(\mult_21_3/ab[1][5] ),
	.B(\mult_21_3/ab[0][6] ),
	.OUT(n213));
   INVERTER U912 (.IN(\mult_21_3/ab[3][4] ),
	.OUT(n1387));
   AOI22 U913 (.A(n1389),
	.B(\mult_21_3/ab[2][4] ),
	.C(n216),
	.D(n852),
	.OUT(n1388));
   INVERTER U914 (.IN(\mult_21_3/ab[4][3] ),
	.OUT(n1390));
   OAI21 U915 (.OUT(n225),
	.C(n1391),
	.B(n1382),
	.A(n1383));
   INVERTER U916 (.IN(\mult_21_3/ab[5][2] ),
	.OUT(n1392));
   OAI21 U917 (.OUT(n233),
	.C(n1393),
	.B(n1392),
	.A(n1385));
   NAND2 U918 (.A(\mult_21_3/ab[1][6] ),
	.B(\mult_21_3/ab[0][7] ),
	.OUT(n1394));
   INVERTER U919 (.IN(\mult_21_3/ab[2][6] ),
	.OUT(n1395));
   INVERTER U920 (.IN(\mult_21_3/ab[1][7] ),
	.OUT(n1396));
   INVERTER U921 (.IN(\mult_21_3/ab[3][5] ),
	.OUT(n1397));
   AOI22 U922 (.A(n1399),
	.B(\mult_21_3/ab[2][5] ),
	.C(n211),
	.D(n851),
	.OUT(n1398));
   INVERTER U923 (.IN(\mult_21_3/ab[4][4] ),
	.OUT(n1400));
   OAI21 U924 (.OUT(n220),
	.C(n1401),
	.B(n1387),
	.A(n1388));
   INVERTER U925 (.IN(\mult_21_3/ab[5][3] ),
	.OUT(n1402));
   OAI22 U926 (.OUT(n1403),
	.D(n865),
	.C(n1390),
	.B(n224),
	.A(n1404));
   OAI22 U927 (.OUT(n235),
	.D(n885),
	.C(n1406),
	.B(n232),
	.A(n1405));
   OAI21 U928 (.OUT(n215),
	.C(n1407),
	.B(n1397),
	.A(n1398));
   INVERTER U929 (.IN(\mult_21_3/ab[5][4] ),
	.OUT(n1408));
   OAI22 U930 (.OUT(n1409),
	.D(n856),
	.C(n1400),
	.B(n219),
	.A(n1410));
   INVERTER U931 (.IN(\mult_21_3/ab[6][3] ),
	.OUT(n1411));
   OAI21 U932 (.OUT(n227),
	.C(n1413),
	.B(n1402),
	.A(n1412));
   INVERTER U933 (.IN(\mult_21_3/ab[5][5] ),
	.OUT(n1414));
   AOI22 U934 (.A(n215),
	.B(\mult_21_3/ab[4][5] ),
	.C(n1416),
	.D(n868),
	.OUT(n1415));
   INVERTER U935 (.IN(\mult_21_3/ab[6][4] ),
	.OUT(n1417));
   OAI21 U936 (.OUT(n264),
	.C(n1419),
	.B(n1408),
	.A(n1418));
   OAI22 U937 (.OUT(n266),
	.D(n871),
	.C(n1411),
	.B(n226),
	.A(n1420));
   NAND2 U938 (.A(\mult_21_3/ab[0][2] ),
	.B(\mult_21_3/ab[1][1] ),
	.OUT(n1421));
   AOI22 U939 (.A(\mult_21_3/ab[2][1] ),
	.B(n237),
	.C(n1423),
	.D(n878),
	.OUT(n1422));
   INVERTER U940 (.IN(\mult_21_3/ab[3][1] ),
	.OUT(n1424));
   OAI21 U941 (.OUT(n239),
	.C(n1425),
	.B(n1424),
	.A(n1422));
   OAI22 U942 (.OUT(n1426),
	.D(n891),
	.C(n1428),
	.B(n238),
	.A(n1427));
   INVERTER U943 (.IN(\mult_21_3/ab[5][1] ),
	.OUT(n1429));
   OAI21 U944 (.OUT(n241),
	.C(n1431),
	.B(n1429),
	.A(n1430));
   OAI22 U945 (.OUT(n243),
	.D(n894),
	.C(n1433),
	.B(n240),
	.A(n1432));
   NAND2 U946 (.A(\mult_21_3/ab[0][1] ),
	.B(\mult_21_3/ab[1][0] ),
	.OUT(n1434));
   AOI22 U947 (.A(\mult_21_3/ab[2][0] ),
	.B(n245),
	.C(n1436),
	.D(n887),
	.OUT(n1435));
   INVERTER U948 (.IN(\mult_21_3/ab[3][0] ),
	.OUT(n1437));
   OAI21 U949 (.OUT(n247),
	.C(n1438),
	.B(n1437),
	.A(n1435));
   INVERTER U950 (.IN(\mult_21_3/ab[4][0] ),
	.OUT(n1439));
   OAI22 U951 (.OUT(n1440),
	.D(n1442),
	.C(n1439),
	.B(n246),
	.A(n1441));
   INVERTER U952 (.IN(\mult_21_3/ab[5][0] ),
	.OUT(n1443));
   OAI21 U953 (.OUT(n249),
	.C(n1445),
	.B(n1443),
	.A(n1444));
   INVERTER U954 (.IN(\mult_21_3/ab[6][0] ),
	.OUT(n1446));
   OAI22 U955 (.OUT(n251),
	.D(n1448),
	.C(n1446),
	.B(n248),
	.A(n1447));
   INVERTER U956 (.IN(\mult_21_3/ab[7][7] ),
	.OUT(n195));
   OAI21 U957 (.OUT(n259),
	.C(n1449),
	.B(n1414),
	.A(n1415));
   AOI22 U958 (.A(n259),
	.B(\mult_21_3/ab[6][5] ),
	.C(n1450),
	.D(n897),
	.OUT(n262));
   INVERTER U959 (.IN(\mult_21_3/ab[7][5] ),
	.OUT(n261));
   OAI22 U960 (.OUT(n1451),
	.D(n873),
	.C(n1417),
	.B(n263),
	.A(n1452));
   INVERTER U961 (.IN(\mult_21_3/ab[7][4] ),
	.OUT(n1453));
   NAND2 U962 (.A(\mult_21_2/ab[0][3] ),
	.B(\mult_21_2/ab[1][2] ),
	.OUT(n1454));
   AOI22 U963 (.A(\mult_21_2/ab[2][2] ),
	.B(n286),
	.C(n1456),
	.D(n918),
	.OUT(n1455));
   NAND2 U964 (.A(\mult_21_2/ab[1][3] ),
	.B(\mult_21_2/ab[0][4] ),
	.OUT(n280));
   INVERTER U965 (.IN(\mult_21_2/ab[3][2] ),
	.OUT(n1457));
   OAI21 U966 (.OUT(n288),
	.C(n1458),
	.B(n1457),
	.A(n1455));
   NAND2 U967 (.A(\mult_21_2/ab[1][4] ),
	.B(\mult_21_2/ab[0][5] ),
	.OUT(n275));
   INVERTER U968 (.IN(\mult_21_2/ab[3][3] ),
	.OUT(n1459));
   AOI22 U969 (.A(n1461),
	.B(\mult_21_2/ab[2][3] ),
	.C(n278),
	.D(n915),
	.OUT(n1460));
   AOI22 U970 (.A(n288),
	.B(\mult_21_2/ab[4][2] ),
	.C(n1463),
	.D(n939),
	.OUT(n1462));
   NAND2 U971 (.A(\mult_21_2/ab[1][5] ),
	.B(\mult_21_2/ab[0][6] ),
	.OUT(n270));
   INVERTER U972 (.IN(\mult_21_2/ab[3][4] ),
	.OUT(n1464));
   AOI22 U973 (.A(n1466),
	.B(\mult_21_2/ab[2][4] ),
	.C(n273),
	.D(n909),
	.OUT(n1465));
   INVERTER U974 (.IN(\mult_21_2/ab[4][3] ),
	.OUT(n1467));
   OAI21 U975 (.OUT(n282),
	.C(n1468),
	.B(n1459),
	.A(n1460));
   INVERTER U976 (.IN(\mult_21_2/ab[5][2] ),
	.OUT(n1469));
   OAI21 U977 (.OUT(n290),
	.C(n1470),
	.B(n1469),
	.A(n1462));
   NAND2 U978 (.A(\mult_21_2/ab[1][6] ),
	.B(\mult_21_2/ab[0][7] ),
	.OUT(n1471));
   INVERTER U979 (.IN(\mult_21_2/ab[2][6] ),
	.OUT(n1472));
   INVERTER U980 (.IN(\mult_21_2/ab[1][7] ),
	.OUT(n1473));
   INVERTER U981 (.IN(\mult_21_2/ab[3][5] ),
	.OUT(n1474));
   AOI22 U982 (.A(n1476),
	.B(\mult_21_2/ab[2][5] ),
	.C(n268),
	.D(n908),
	.OUT(n1475));
   INVERTER U983 (.IN(\mult_21_2/ab[4][4] ),
	.OUT(n1477));
   OAI21 U984 (.OUT(n277),
	.C(n1478),
	.B(n1464),
	.A(n1465));
   INVERTER U985 (.IN(\mult_21_2/ab[5][3] ),
	.OUT(n1479));
   OAI22 U986 (.OUT(n1480),
	.D(n922),
	.C(n1467),
	.B(n281),
	.A(n1481));
   OAI22 U987 (.OUT(n292),
	.D(n942),
	.C(n1483),
	.B(n289),
	.A(n1482));
   OAI21 U988 (.OUT(n272),
	.C(n1484),
	.B(n1474),
	.A(n1475));
   INVERTER U989 (.IN(\mult_21_2/ab[5][4] ),
	.OUT(n1485));
   OAI22 U990 (.OUT(n1486),
	.D(n913),
	.C(n1477),
	.B(n276),
	.A(n1487));
   INVERTER U991 (.IN(\mult_21_2/ab[6][3] ),
	.OUT(n1488));
   OAI21 U992 (.OUT(n284),
	.C(n1490),
	.B(n1479),
	.A(n1489));
   INVERTER U993 (.IN(\mult_21_2/ab[5][5] ),
	.OUT(n1491));
   AOI22 U994 (.A(n272),
	.B(\mult_21_2/ab[4][5] ),
	.C(n1493),
	.D(n925),
	.OUT(n1492));
   INVERTER U995 (.IN(\mult_21_2/ab[6][4] ),
	.OUT(n1494));
   OAI21 U996 (.OUT(n321),
	.C(n1496),
	.B(n1485),
	.A(n1495));
   OAI22 U997 (.OUT(n323),
	.D(n928),
	.C(n1488),
	.B(n283),
	.A(n1497));
   NAND2 U998 (.A(\mult_21_2/ab[0][2] ),
	.B(\mult_21_2/ab[1][1] ),
	.OUT(n1498));
   AOI22 U999 (.A(\mult_21_2/ab[2][1] ),
	.B(n294),
	.C(n1500),
	.D(n935),
	.OUT(n1499));
   INVERTER U1000 (.IN(\mult_21_2/ab[3][1] ),
	.OUT(n1501));
   OAI21 U1001 (.OUT(n296),
	.C(n1502),
	.B(n1501),
	.A(n1499));
   OAI22 U1002 (.OUT(n1503),
	.D(n948),
	.C(n1505),
	.B(n295),
	.A(n1504));
   INVERTER U1003 (.IN(\mult_21_2/ab[5][1] ),
	.OUT(n1506));
   OAI21 U1004 (.OUT(n298),
	.C(n1508),
	.B(n1506),
	.A(n1507));
   OAI22 U1005 (.OUT(n300),
	.D(n951),
	.C(n1510),
	.B(n297),
	.A(n1509));
   NAND2 U1006 (.A(\mult_21_2/ab[0][1] ),
	.B(\mult_21_2/ab[1][0] ),
	.OUT(n1511));
   AOI22 U1007 (.A(\mult_21_2/ab[2][0] ),
	.B(n302),
	.C(n1513),
	.D(n944),
	.OUT(n1512));
   INVERTER U1008 (.IN(\mult_21_2/ab[3][0] ),
	.OUT(n1514));
   OAI21 U1009 (.OUT(n304),
	.C(n1515),
	.B(n1514),
	.A(n1512));
   INVERTER U1010 (.IN(\mult_21_2/ab[4][0] ),
	.OUT(n1516));
   OAI22 U1011 (.OUT(n1517),
	.D(n1519),
	.C(n1516),
	.B(n303),
	.A(n1518));
   INVERTER U1012 (.IN(\mult_21_2/ab[5][0] ),
	.OUT(n1520));
   OAI21 U1013 (.OUT(n306),
	.C(n1522),
	.B(n1520),
	.A(n1521));
   INVERTER U1014 (.IN(\mult_21_2/ab[6][0] ),
	.OUT(n1523));
   OAI22 U1015 (.OUT(n308),
	.D(n1525),
	.C(n1523),
	.B(n305),
	.A(n1524));
   INVERTER U1016 (.IN(\mult_21_2/ab[7][7] ),
	.OUT(n179));
   OAI21 U1017 (.OUT(n316),
	.C(n1526),
	.B(n1491),
	.A(n1492));
   AOI22 U1018 (.A(n316),
	.B(\mult_21_2/ab[6][5] ),
	.C(n1527),
	.D(n954),
	.OUT(n319));
   INVERTER U1019 (.IN(\mult_21_2/ab[7][5] ),
	.OUT(n318));
   OAI22 U1020 (.OUT(n1528),
	.D(n930),
	.C(n1494),
	.B(n320),
	.A(n1529));
   INVERTER U1021 (.IN(\mult_21_2/ab[7][4] ),
	.OUT(n1530));
   NAND2 U1022 (.A(\mult_21/ab[0][3] ),
	.B(\mult_21/ab[1][2] ),
	.OUT(n1531));
   AOI22 U1023 (.A(\mult_21/ab[2][2] ),
	.B(n343),
	.C(n1533),
	.D(n975),
	.OUT(n1532));
   NAND2 U1024 (.A(\mult_21/ab[1][3] ),
	.B(\mult_21/ab[0][4] ),
	.OUT(n337));
   INVERTER U1025 (.IN(\mult_21/ab[3][2] ),
	.OUT(n1534));
   OAI21 U1026 (.OUT(n345),
	.C(n1535),
	.B(n1534),
	.A(n1532));
   NAND2 U1027 (.A(\mult_21/ab[1][4] ),
	.B(\mult_21/ab[0][5] ),
	.OUT(n332));
   INVERTER U1028 (.IN(\mult_21/ab[3][3] ),
	.OUT(n1536));
   AOI22 U1029 (.A(n1538),
	.B(\mult_21/ab[2][3] ),
	.C(n335),
	.D(n972),
	.OUT(n1537));
   AOI22 U1030 (.A(n345),
	.B(\mult_21/ab[4][2] ),
	.C(n1540),
	.D(n996),
	.OUT(n1539));
   NAND2 U1031 (.A(\mult_21/ab[1][5] ),
	.B(\mult_21/ab[0][6] ),
	.OUT(n327));
   INVERTER U1032 (.IN(\mult_21/ab[3][4] ),
	.OUT(n1541));
   AOI22 U1033 (.A(n1543),
	.B(\mult_21/ab[2][4] ),
	.C(n330),
	.D(n966),
	.OUT(n1542));
   INVERTER U1034 (.IN(\mult_21/ab[4][3] ),
	.OUT(n1544));
   OAI21 U1035 (.OUT(n339),
	.C(n1545),
	.B(n1536),
	.A(n1537));
   INVERTER U1036 (.IN(\mult_21/ab[5][2] ),
	.OUT(n1546));
   OAI21 U1037 (.OUT(n347),
	.C(n1547),
	.B(n1546),
	.A(n1539));
   NAND2 U1038 (.A(\mult_21/ab[1][6] ),
	.B(\mult_21/ab[0][7] ),
	.OUT(n1548));
   INVERTER U1039 (.IN(\mult_21/ab[2][6] ),
	.OUT(n1549));
   INVERTER U1040 (.IN(\mult_21/ab[1][7] ),
	.OUT(n1550));
   INVERTER U1041 (.IN(\mult_21/ab[3][5] ),
	.OUT(n1551));
   AOI22 U1042 (.A(n1553),
	.B(\mult_21/ab[2][5] ),
	.C(n325),
	.D(n965),
	.OUT(n1552));
   INVERTER U1043 (.IN(\mult_21/ab[4][4] ),
	.OUT(n1554));
   OAI21 U1044 (.OUT(n334),
	.C(n1555),
	.B(n1541),
	.A(n1542));
   INVERTER U1045 (.IN(\mult_21/ab[5][3] ),
	.OUT(n1556));
   OAI22 U1046 (.OUT(n1557),
	.D(n979),
	.C(n1544),
	.B(n338),
	.A(n1558));
   OAI22 U1047 (.OUT(n349),
	.D(n999),
	.C(n1560),
	.B(n346),
	.A(n1559));
   OAI21 U1048 (.OUT(n329),
	.C(n1561),
	.B(n1551),
	.A(n1552));
   INVERTER U1049 (.IN(\mult_21/ab[5][4] ),
	.OUT(n1562));
   OAI22 U1050 (.OUT(n1563),
	.D(n970),
	.C(n1554),
	.B(n333),
	.A(n1564));
   INVERTER U1051 (.IN(\mult_21/ab[6][3] ),
	.OUT(n1565));
   OAI21 U1052 (.OUT(n341),
	.C(n1567),
	.B(n1556),
	.A(n1566));
   INVERTER U1053 (.IN(\mult_21/ab[5][5] ),
	.OUT(n1568));
   AOI22 U1054 (.A(n329),
	.B(\mult_21/ab[4][5] ),
	.C(n1570),
	.D(n982),
	.OUT(n1569));
   INVERTER U1055 (.IN(\mult_21/ab[6][4] ),
	.OUT(n1571));
   OAI21 U1056 (.OUT(n378),
	.C(n1573),
	.B(n1562),
	.A(n1572));
   OAI22 U1057 (.OUT(n380),
	.D(n985),
	.C(n1565),
	.B(n340),
	.A(n1574));
   NAND2 U1058 (.A(\mult_21/ab[0][2] ),
	.B(\mult_21/ab[1][1] ),
	.OUT(n1575));
   AOI22 U1059 (.A(\mult_21/ab[2][1] ),
	.B(n351),
	.C(n1577),
	.D(n992),
	.OUT(n1576));
   INVERTER U1060 (.IN(\mult_21/ab[3][1] ),
	.OUT(n1578));
   OAI21 U1061 (.OUT(n353),
	.C(n1579),
	.B(n1578),
	.A(n1576));
   OAI22 U1062 (.OUT(n1580),
	.D(n1005),
	.C(n1582),
	.B(n352),
	.A(n1581));
   INVERTER U1063 (.IN(\mult_21/ab[5][1] ),
	.OUT(n1583));
   OAI21 U1064 (.OUT(n355),
	.C(n1585),
	.B(n1583),
	.A(n1584));
   OAI22 U1065 (.OUT(n357),
	.D(n1008),
	.C(n1587),
	.B(n354),
	.A(n1586));
   NAND2 U1066 (.A(\mult_21/ab[0][1] ),
	.B(\mult_21/ab[1][0] ),
	.OUT(n1588));
   AOI22 U1067 (.A(\mult_21/ab[2][0] ),
	.B(n359),
	.C(n1590),
	.D(n1001),
	.OUT(n1589));
   INVERTER U1068 (.IN(\mult_21/ab[3][0] ),
	.OUT(n1591));
   OAI21 U1069 (.OUT(n361),
	.C(n1592),
	.B(n1591),
	.A(n1589));
   INVERTER U1070 (.IN(\mult_21/ab[4][0] ),
	.OUT(n1593));
   OAI22 U1071 (.OUT(n1594),
	.D(n1596),
	.C(n1593),
	.B(n360),
	.A(n1595));
   INVERTER U1072 (.IN(\mult_21/ab[5][0] ),
	.OUT(n1597));
   OAI21 U1073 (.OUT(n363),
	.C(n1599),
	.B(n1597),
	.A(n1598));
   INVERTER U1074 (.IN(\mult_21/ab[6][0] ),
	.OUT(n1600));
   OAI22 U1075 (.OUT(n365),
	.D(n1602),
	.C(n1600),
	.B(n362),
	.A(n1601));
   INVERTER U1076 (.IN(\mult_21/ab[7][7] ),
	.OUT(n163));
   OAI21 U1077 (.OUT(n373),
	.C(n1603),
	.B(n1568),
	.A(n1569));
   AOI22 U1078 (.A(n373),
	.B(\mult_21/ab[6][5] ),
	.C(n1604),
	.D(n1011),
	.OUT(n376));
   INVERTER U1079 (.IN(\mult_21/ab[7][5] ),
	.OUT(n375));
   OAI22 U1080 (.OUT(n1605),
	.D(n987),
	.C(n1571),
	.B(n377),
	.A(n1606));
   INVERTER U1081 (.IN(\mult_21/ab[7][4] ),
	.OUT(n1607));
   NAND2 U1082 (.A(\mult_20_3/ab[0][3] ),
	.B(\mult_20_3/ab[1][2] ),
	.OUT(n1608));
   AOI22 U1083 (.A(\mult_20_3/ab[2][2] ),
	.B(n400),
	.C(n1610),
	.D(n1032),
	.OUT(n1609));
   NAND2 U1084 (.A(\mult_20_3/ab[1][3] ),
	.B(\mult_20_3/ab[0][4] ),
	.OUT(n394));
   INVERTER U1085 (.IN(\mult_20_3/ab[3][2] ),
	.OUT(n1611));
   OAI21 U1086 (.OUT(n402),
	.C(n1612),
	.B(n1611),
	.A(n1609));
   NAND2 U1087 (.A(\mult_20_3/ab[1][4] ),
	.B(\mult_20_3/ab[0][5] ),
	.OUT(n389));
   INVERTER U1088 (.IN(\mult_20_3/ab[3][3] ),
	.OUT(n1613));
   AOI22 U1089 (.A(n1615),
	.B(\mult_20_3/ab[2][3] ),
	.C(n392),
	.D(n1029),
	.OUT(n1614));
   AOI22 U1090 (.A(n402),
	.B(\mult_20_3/ab[4][2] ),
	.C(n1617),
	.D(n1053),
	.OUT(n1616));
   NAND2 U1091 (.A(\mult_20_3/ab[1][5] ),
	.B(\mult_20_3/ab[0][6] ),
	.OUT(n384));
   INVERTER U1092 (.IN(\mult_20_3/ab[3][4] ),
	.OUT(n1618));
   AOI22 U1093 (.A(n1620),
	.B(\mult_20_3/ab[2][4] ),
	.C(n387),
	.D(n1023),
	.OUT(n1619));
   INVERTER U1094 (.IN(\mult_20_3/ab[4][3] ),
	.OUT(n1621));
   OAI21 U1095 (.OUT(n396),
	.C(n1622),
	.B(n1613),
	.A(n1614));
   INVERTER U1096 (.IN(\mult_20_3/ab[5][2] ),
	.OUT(n1623));
   OAI21 U1097 (.OUT(n404),
	.C(n1624),
	.B(n1623),
	.A(n1616));
   NAND2 U1098 (.A(\mult_20_3/ab[1][6] ),
	.B(\mult_20_3/ab[0][7] ),
	.OUT(n1625));
   INVERTER U1099 (.IN(\mult_20_3/ab[2][6] ),
	.OUT(n1626));
   INVERTER U1100 (.IN(\mult_20_3/ab[1][7] ),
	.OUT(n1627));
   INVERTER U1101 (.IN(\mult_20_3/ab[3][5] ),
	.OUT(n1628));
   AOI22 U1102 (.A(n1630),
	.B(\mult_20_3/ab[2][5] ),
	.C(n382),
	.D(n1022),
	.OUT(n1629));
   INVERTER U1103 (.IN(\mult_20_3/ab[4][4] ),
	.OUT(n1631));
   OAI21 U1104 (.OUT(n391),
	.C(n1632),
	.B(n1618),
	.A(n1619));
   INVERTER U1105 (.IN(\mult_20_3/ab[5][3] ),
	.OUT(n1633));
   OAI22 U1106 (.OUT(n1634),
	.D(n1036),
	.C(n1621),
	.B(n395),
	.A(n1635));
   OAI22 U1107 (.OUT(n406),
	.D(n1056),
	.C(n1637),
	.B(n403),
	.A(n1636));
   OAI21 U1108 (.OUT(n386),
	.C(n1638),
	.B(n1628),
	.A(n1629));
   INVERTER U1109 (.IN(\mult_20_3/ab[5][4] ),
	.OUT(n1639));
   OAI22 U1110 (.OUT(n1640),
	.D(n1027),
	.C(n1631),
	.B(n390),
	.A(n1641));
   INVERTER U1111 (.IN(\mult_20_3/ab[6][3] ),
	.OUT(n1642));
   OAI21 U1112 (.OUT(n398),
	.C(n1644),
	.B(n1633),
	.A(n1643));
   INVERTER U1113 (.IN(\mult_20_3/ab[5][5] ),
	.OUT(n1645));
   AOI22 U1114 (.A(n386),
	.B(\mult_20_3/ab[4][5] ),
	.C(n1647),
	.D(n1039),
	.OUT(n1646));
   INVERTER U1115 (.IN(\mult_20_3/ab[6][4] ),
	.OUT(n1648));
   OAI21 U1116 (.OUT(n435),
	.C(n1650),
	.B(n1639),
	.A(n1649));
   OAI22 U1117 (.OUT(n437),
	.D(n1042),
	.C(n1642),
	.B(n397),
	.A(n1651));
   NAND2 U1118 (.A(\mult_20_3/ab[0][2] ),
	.B(\mult_20_3/ab[1][1] ),
	.OUT(n1652));
   AOI22 U1119 (.A(\mult_20_3/ab[2][1] ),
	.B(n408),
	.C(n1654),
	.D(n1049),
	.OUT(n1653));
   INVERTER U1120 (.IN(\mult_20_3/ab[3][1] ),
	.OUT(n1655));
   OAI21 U1121 (.OUT(n410),
	.C(n1656),
	.B(n1655),
	.A(n1653));
   OAI22 U1122 (.OUT(n1657),
	.D(n1062),
	.C(n1659),
	.B(n409),
	.A(n1658));
   INVERTER U1123 (.IN(\mult_20_3/ab[5][1] ),
	.OUT(n1660));
   OAI21 U1124 (.OUT(n412),
	.C(n1662),
	.B(n1660),
	.A(n1661));
   OAI22 U1125 (.OUT(n414),
	.D(n1065),
	.C(n1664),
	.B(n411),
	.A(n1663));
   NAND2 U1126 (.A(\mult_20_3/ab[0][1] ),
	.B(\mult_20_3/ab[1][0] ),
	.OUT(n1665));
   AOI22 U1127 (.A(\mult_20_3/ab[2][0] ),
	.B(n416),
	.C(n1667),
	.D(n1058),
	.OUT(n1666));
   INVERTER U1128 (.IN(\mult_20_3/ab[3][0] ),
	.OUT(n1668));
   OAI21 U1129 (.OUT(n418),
	.C(n1669),
	.B(n1668),
	.A(n1666));
   INVERTER U1130 (.IN(\mult_20_3/ab[4][0] ),
	.OUT(n1670));
   OAI22 U1131 (.OUT(n1671),
	.D(n1673),
	.C(n1670),
	.B(n417),
	.A(n1672));
   INVERTER U1132 (.IN(\mult_20_3/ab[5][0] ),
	.OUT(n1674));
   OAI21 U1133 (.OUT(n420),
	.C(n1676),
	.B(n1674),
	.A(n1675));
   INVERTER U1134 (.IN(\mult_20_3/ab[6][0] ),
	.OUT(n1677));
   OAI22 U1135 (.OUT(n422),
	.D(n1679),
	.C(n1677),
	.B(n419),
	.A(n1678));
   INVERTER U1136 (.IN(\mult_20_3/ab[7][7] ),
	.OUT(n147));
   OAI21 U1137 (.OUT(n430),
	.C(n1680),
	.B(n1645),
	.A(n1646));
   AOI22 U1138 (.A(n430),
	.B(\mult_20_3/ab[6][5] ),
	.C(n1681),
	.D(n1068),
	.OUT(n433));
   INVERTER U1139 (.IN(\mult_20_3/ab[7][5] ),
	.OUT(n432));
   OAI22 U1140 (.OUT(n1682),
	.D(n1044),
	.C(n1648),
	.B(n434),
	.A(n1683));
   INVERTER U1141 (.IN(\mult_20_3/ab[7][4] ),
	.OUT(n1684));
   NAND2 U1142 (.A(\mult_20_2/ab[0][3] ),
	.B(\mult_20_2/ab[1][2] ),
	.OUT(n1685));
   AOI22 U1143 (.A(\mult_20_2/ab[2][2] ),
	.B(n457),
	.C(n1687),
	.D(n1089),
	.OUT(n1686));
   NAND2 U1144 (.A(\mult_20_2/ab[1][3] ),
	.B(\mult_20_2/ab[0][4] ),
	.OUT(n451));
   INVERTER U1145 (.IN(\mult_20_2/ab[3][2] ),
	.OUT(n1688));
   OAI21 U1146 (.OUT(n459),
	.C(n1689),
	.B(n1688),
	.A(n1686));
   NAND2 U1147 (.A(\mult_20_2/ab[1][4] ),
	.B(\mult_20_2/ab[0][5] ),
	.OUT(n446));
   INVERTER U1148 (.IN(\mult_20_2/ab[3][3] ),
	.OUT(n1690));
   AOI22 U1149 (.A(n1692),
	.B(\mult_20_2/ab[2][3] ),
	.C(n449),
	.D(n1086),
	.OUT(n1691));
   AOI22 U1150 (.A(n459),
	.B(\mult_20_2/ab[4][2] ),
	.C(n1694),
	.D(n1110),
	.OUT(n1693));
   NAND2 U1151 (.A(\mult_20_2/ab[1][5] ),
	.B(\mult_20_2/ab[0][6] ),
	.OUT(n441));
   INVERTER U1152 (.IN(\mult_20_2/ab[3][4] ),
	.OUT(n1695));
   AOI22 U1153 (.A(n1697),
	.B(\mult_20_2/ab[2][4] ),
	.C(n444),
	.D(n1080),
	.OUT(n1696));
   INVERTER U1154 (.IN(\mult_20_2/ab[4][3] ),
	.OUT(n1698));
   OAI21 U1155 (.OUT(n453),
	.C(n1699),
	.B(n1690),
	.A(n1691));
   INVERTER U1156 (.IN(\mult_20_2/ab[5][2] ),
	.OUT(n1700));
   OAI21 U1157 (.OUT(n461),
	.C(n1701),
	.B(n1700),
	.A(n1693));
   NAND2 U1158 (.A(\mult_20_2/ab[1][6] ),
	.B(\mult_20_2/ab[0][7] ),
	.OUT(n1702));
   INVERTER U1159 (.IN(\mult_20_2/ab[2][6] ),
	.OUT(n1703));
   INVERTER U1160 (.IN(\mult_20_2/ab[1][7] ),
	.OUT(n1704));
   INVERTER U1161 (.IN(\mult_20_2/ab[3][5] ),
	.OUT(n1705));
   AOI22 U1162 (.A(n1707),
	.B(\mult_20_2/ab[2][5] ),
	.C(n439),
	.D(n1079),
	.OUT(n1706));
   INVERTER U1163 (.IN(\mult_20_2/ab[4][4] ),
	.OUT(n1708));
   OAI21 U1164 (.OUT(n448),
	.C(n1709),
	.B(n1695),
	.A(n1696));
   INVERTER U1165 (.IN(\mult_20_2/ab[5][3] ),
	.OUT(n1710));
   OAI22 U1166 (.OUT(n1711),
	.D(n1093),
	.C(n1698),
	.B(n452),
	.A(n1712));
   OAI22 U1167 (.OUT(n463),
	.D(n1113),
	.C(n1714),
	.B(n460),
	.A(n1713));
   OAI21 U1168 (.OUT(n443),
	.C(n1715),
	.B(n1705),
	.A(n1706));
   INVERTER U1169 (.IN(\mult_20_2/ab[5][4] ),
	.OUT(n1716));
   OAI22 U1170 (.OUT(n1717),
	.D(n1084),
	.C(n1708),
	.B(n447),
	.A(n1718));
   INVERTER U1171 (.IN(\mult_20_2/ab[6][3] ),
	.OUT(n1719));
   OAI21 U1172 (.OUT(n455),
	.C(n1721),
	.B(n1710),
	.A(n1720));
   INVERTER U1173 (.IN(\mult_20_2/ab[5][5] ),
	.OUT(n1722));
   AOI22 U1174 (.A(n443),
	.B(\mult_20_2/ab[4][5] ),
	.C(n1724),
	.D(n1096),
	.OUT(n1723));
   INVERTER U1175 (.IN(\mult_20_2/ab[6][4] ),
	.OUT(n1725));
   OAI21 U1176 (.OUT(n492),
	.C(n1727),
	.B(n1716),
	.A(n1726));
   OAI22 U1177 (.OUT(n494),
	.D(n1099),
	.C(n1719),
	.B(n454),
	.A(n1728));
   NAND2 U1178 (.A(\mult_20_2/ab[0][2] ),
	.B(\mult_20_2/ab[1][1] ),
	.OUT(n1729));
   AOI22 U1179 (.A(\mult_20_2/ab[2][1] ),
	.B(n465),
	.C(n1731),
	.D(n1106),
	.OUT(n1730));
   INVERTER U1180 (.IN(\mult_20_2/ab[3][1] ),
	.OUT(n1732));
   OAI21 U1181 (.OUT(n467),
	.C(n1733),
	.B(n1732),
	.A(n1730));
   OAI22 U1182 (.OUT(n1734),
	.D(n1119),
	.C(n1736),
	.B(n466),
	.A(n1735));
   INVERTER U1183 (.IN(\mult_20_2/ab[5][1] ),
	.OUT(n1737));
   OAI21 U1184 (.OUT(n469),
	.C(n1739),
	.B(n1737),
	.A(n1738));
   OAI22 U1185 (.OUT(n471),
	.D(n1122),
	.C(n1741),
	.B(n468),
	.A(n1740));
   NAND2 U1186 (.A(\mult_20_2/ab[0][1] ),
	.B(\mult_20_2/ab[1][0] ),
	.OUT(n1742));
   AOI22 U1187 (.A(\mult_20_2/ab[2][0] ),
	.B(n473),
	.C(n1744),
	.D(n1115),
	.OUT(n1743));
   INVERTER U1188 (.IN(\mult_20_2/ab[3][0] ),
	.OUT(n1745));
   OAI21 U1189 (.OUT(n475),
	.C(n1746),
	.B(n1745),
	.A(n1743));
   INVERTER U1190 (.IN(\mult_20_2/ab[4][0] ),
	.OUT(n1747));
   OAI22 U1191 (.OUT(n1748),
	.D(n1750),
	.C(n1747),
	.B(n474),
	.A(n1749));
   INVERTER U1192 (.IN(\mult_20_2/ab[5][0] ),
	.OUT(n1751));
   OAI21 U1193 (.OUT(n477),
	.C(n1753),
	.B(n1751),
	.A(n1752));
   INVERTER U1194 (.IN(\mult_20_2/ab[6][0] ),
	.OUT(n1754));
   OAI22 U1195 (.OUT(n479),
	.D(n1756),
	.C(n1754),
	.B(n476),
	.A(n1755));
   INVERTER U1196 (.IN(\mult_20_2/ab[7][7] ),
	.OUT(n131));
   OAI21 U1197 (.OUT(n487),
	.C(n1757),
	.B(n1722),
	.A(n1723));
   AOI22 U1198 (.A(n487),
	.B(\mult_20_2/ab[6][5] ),
	.C(n1758),
	.D(n1125),
	.OUT(n490));
   INVERTER U1199 (.IN(\mult_20_2/ab[7][5] ),
	.OUT(n489));
   OAI22 U1200 (.OUT(n1759),
	.D(n1101),
	.C(n1725),
	.B(n491),
	.A(n1760));
   INVERTER U1201 (.IN(\mult_20_2/ab[7][4] ),
	.OUT(n1761));
   NAND2 U1202 (.A(\mult_20/ab[0][3] ),
	.B(\mult_20/ab[1][2] ),
	.OUT(n1762));
   AOI22 U1203 (.A(\mult_20/ab[2][2] ),
	.B(n514),
	.C(n1764),
	.D(n1146),
	.OUT(n1763));
   NAND2 U1204 (.A(\mult_20/ab[1][3] ),
	.B(\mult_20/ab[0][4] ),
	.OUT(n508));
   INVERTER U1205 (.IN(\mult_20/ab[3][2] ),
	.OUT(n1765));
   OAI21 U1206 (.OUT(n516),
	.C(n1766),
	.B(n1765),
	.A(n1763));
   NAND2 U1207 (.A(\mult_20/ab[1][4] ),
	.B(\mult_20/ab[0][5] ),
	.OUT(n503));
   INVERTER U1208 (.IN(\mult_20/ab[3][3] ),
	.OUT(n1767));
   AOI22 U1209 (.A(n1769),
	.B(\mult_20/ab[2][3] ),
	.C(n506),
	.D(n1143),
	.OUT(n1768));
   AOI22 U1210 (.A(n516),
	.B(\mult_20/ab[4][2] ),
	.C(n1771),
	.D(n1167),
	.OUT(n1770));
   NAND2 U1211 (.A(\mult_20/ab[1][5] ),
	.B(\mult_20/ab[0][6] ),
	.OUT(n498));
   INVERTER U1212 (.IN(\mult_20/ab[3][4] ),
	.OUT(n1772));
   AOI22 U1213 (.A(n1774),
	.B(\mult_20/ab[2][4] ),
	.C(n501),
	.D(n1137),
	.OUT(n1773));
   INVERTER U1214 (.IN(\mult_20/ab[4][3] ),
	.OUT(n1775));
   OAI21 U1215 (.OUT(n510),
	.C(n1776),
	.B(n1767),
	.A(n1768));
   INVERTER U1216 (.IN(\mult_20/ab[5][2] ),
	.OUT(n1777));
   OAI21 U1217 (.OUT(n518),
	.C(n1778),
	.B(n1777),
	.A(n1770));
   NAND2 U1218 (.A(\mult_20/ab[1][6] ),
	.B(\mult_20/ab[0][7] ),
	.OUT(n1779));
   INVERTER U1219 (.IN(\mult_20/ab[2][6] ),
	.OUT(n1780));
   INVERTER U1220 (.IN(\mult_20/ab[1][7] ),
	.OUT(n1781));
   INVERTER U1221 (.IN(\mult_20/ab[3][5] ),
	.OUT(n1782));
   AOI22 U1222 (.A(n1784),
	.B(\mult_20/ab[2][5] ),
	.C(n496),
	.D(n1136),
	.OUT(n1783));
   INVERTER U1223 (.IN(\mult_20/ab[4][4] ),
	.OUT(n1785));
   OAI21 U1224 (.OUT(n505),
	.C(n1786),
	.B(n1772),
	.A(n1773));
   INVERTER U1225 (.IN(\mult_20/ab[5][3] ),
	.OUT(n1787));
   OAI22 U1226 (.OUT(n1788),
	.D(n1150),
	.C(n1775),
	.B(n509),
	.A(n1789));
   OAI22 U1227 (.OUT(n520),
	.D(n1170),
	.C(n1791),
	.B(n517),
	.A(n1790));
   OAI21 U1228 (.OUT(n500),
	.C(n1792),
	.B(n1782),
	.A(n1783));
   INVERTER U1229 (.IN(\mult_20/ab[5][4] ),
	.OUT(n1793));
   OAI22 U1230 (.OUT(n1794),
	.D(n1141),
	.C(n1785),
	.B(n504),
	.A(n1795));
   INVERTER U1231 (.IN(\mult_20/ab[6][3] ),
	.OUT(n1796));
   OAI21 U1232 (.OUT(n512),
	.C(n1798),
	.B(n1787),
	.A(n1797));
   INVERTER U1233 (.IN(\mult_20/ab[5][5] ),
	.OUT(n1799));
   AOI22 U1234 (.A(n500),
	.B(\mult_20/ab[4][5] ),
	.C(n1801),
	.D(n1153),
	.OUT(n1800));
   INVERTER U1235 (.IN(\mult_20/ab[6][4] ),
	.OUT(n1802));
   OAI21 U1236 (.OUT(n549),
	.C(n1804),
	.B(n1793),
	.A(n1803));
   OAI22 U1237 (.OUT(n551),
	.D(n1156),
	.C(n1796),
	.B(n511),
	.A(n1805));
   NAND2 U1238 (.A(\mult_20/ab[0][2] ),
	.B(\mult_20/ab[1][1] ),
	.OUT(n1806));
   AOI22 U1239 (.A(\mult_20/ab[2][1] ),
	.B(n522),
	.C(n1808),
	.D(n1163),
	.OUT(n1807));
   INVERTER U1240 (.IN(\mult_20/ab[3][1] ),
	.OUT(n1809));
   OAI21 U1241 (.OUT(n524),
	.C(n1810),
	.B(n1809),
	.A(n1807));
   OAI22 U1242 (.OUT(n1811),
	.D(n1176),
	.C(n1813),
	.B(n523),
	.A(n1812));
   INVERTER U1243 (.IN(\mult_20/ab[5][1] ),
	.OUT(n1814));
   OAI21 U1244 (.OUT(n526),
	.C(n1816),
	.B(n1814),
	.A(n1815));
   OAI22 U1245 (.OUT(n528),
	.D(n1179),
	.C(n1818),
	.B(n525),
	.A(n1817));
   NAND2 U1246 (.A(\mult_20/ab[0][1] ),
	.B(\mult_20/ab[1][0] ),
	.OUT(n1819));
   AOI22 U1247 (.A(\mult_20/ab[2][0] ),
	.B(n530),
	.C(n1821),
	.D(n1172),
	.OUT(n1820));
   INVERTER U1248 (.IN(\mult_20/ab[3][0] ),
	.OUT(n1822));
   OAI21 U1249 (.OUT(n532),
	.C(n1823),
	.B(n1822),
	.A(n1820));
   INVERTER U1250 (.IN(\mult_20/ab[4][0] ),
	.OUT(n1824));
   OAI22 U1251 (.OUT(n1825),
	.D(n1827),
	.C(n1824),
	.B(n531),
	.A(n1826));
   INVERTER U1252 (.IN(\mult_20/ab[5][0] ),
	.OUT(n1828));
   OAI21 U1253 (.OUT(n534),
	.C(n1830),
	.B(n1828),
	.A(n1829));
   INVERTER U1254 (.IN(\mult_20/ab[6][0] ),
	.OUT(n1831));
   OAI22 U1255 (.OUT(n536),
	.D(n1833),
	.C(n1831),
	.B(n533),
	.A(n1832));
   INVERTER U1256 (.IN(\mult_20/ab[7][7] ),
	.OUT(n115));
   OAI21 U1257 (.OUT(n544),
	.C(n1834),
	.B(n1799),
	.A(n1800));
   AOI22 U1258 (.A(n544),
	.B(\mult_20/ab[6][5] ),
	.C(n1835),
	.D(n1182),
	.OUT(n547));
   INVERTER U1259 (.IN(\mult_20/ab[7][5] ),
	.OUT(n546));
   OAI22 U1260 (.OUT(n1836),
	.D(n1158),
	.C(n1802),
	.B(n548),
	.A(n1837));
   INVERTER U1261 (.IN(\mult_20/ab[7][4] ),
	.OUT(n1838));
   NAND2 U1262 (.A(\mult_19_3/ab[0][3] ),
	.B(\mult_19_3/ab[1][2] ),
	.OUT(n1839));
   AOI22 U1263 (.A(\mult_19_3/ab[2][2] ),
	.B(n571),
	.C(n1841),
	.D(n1203),
	.OUT(n1840));
   NAND2 U1264 (.A(\mult_19_3/ab[1][3] ),
	.B(\mult_19_3/ab[0][4] ),
	.OUT(n565));
   INVERTER U1265 (.IN(\mult_19_3/ab[3][2] ),
	.OUT(n1842));
   OAI21 U1266 (.OUT(n573),
	.C(n1843),
	.B(n1842),
	.A(n1840));
   NAND2 U1267 (.A(\mult_19_3/ab[1][4] ),
	.B(\mult_19_3/ab[0][5] ),
	.OUT(n560));
   INVERTER U1268 (.IN(\mult_19_3/ab[3][3] ),
	.OUT(n1844));
   AOI22 U1269 (.A(n1846),
	.B(\mult_19_3/ab[2][3] ),
	.C(n563),
	.D(n1200),
	.OUT(n1845));
   AOI22 U1270 (.A(n573),
	.B(\mult_19_3/ab[4][2] ),
	.C(n1848),
	.D(n1224),
	.OUT(n1847));
   NAND2 U1271 (.A(\mult_19_3/ab[1][5] ),
	.B(\mult_19_3/ab[0][6] ),
	.OUT(n555));
   INVERTER U1272 (.IN(\mult_19_3/ab[3][4] ),
	.OUT(n1849));
   AOI22 U1273 (.A(n1851),
	.B(\mult_19_3/ab[2][4] ),
	.C(n558),
	.D(n1194),
	.OUT(n1850));
   INVERTER U1274 (.IN(\mult_19_3/ab[4][3] ),
	.OUT(n1852));
   OAI21 U1275 (.OUT(n567),
	.C(n1853),
	.B(n1844),
	.A(n1845));
   INVERTER U1276 (.IN(\mult_19_3/ab[5][2] ),
	.OUT(n1854));
   OAI21 U1277 (.OUT(n575),
	.C(n1855),
	.B(n1854),
	.A(n1847));
   NAND2 U1278 (.A(\mult_19_3/ab[1][6] ),
	.B(\mult_19_3/ab[0][7] ),
	.OUT(n1856));
   INVERTER U1279 (.IN(\mult_19_3/ab[2][6] ),
	.OUT(n1857));
   INVERTER U1280 (.IN(\mult_19_3/ab[1][7] ),
	.OUT(n1858));
   INVERTER U1281 (.IN(\mult_19_3/ab[3][5] ),
	.OUT(n1859));
   AOI22 U1282 (.A(n1861),
	.B(\mult_19_3/ab[2][5] ),
	.C(n553),
	.D(n1193),
	.OUT(n1860));
   INVERTER U1283 (.IN(\mult_19_3/ab[4][4] ),
	.OUT(n1862));
   OAI21 U1284 (.OUT(n562),
	.C(n1863),
	.B(n1849),
	.A(n1850));
   INVERTER U1285 (.IN(\mult_19_3/ab[5][3] ),
	.OUT(n1864));
   OAI22 U1286 (.OUT(n1865),
	.D(n1207),
	.C(n1852),
	.B(n566),
	.A(n1866));
   OAI22 U1287 (.OUT(n577),
	.D(n1227),
	.C(n1868),
	.B(n574),
	.A(n1867));
   OAI21 U1288 (.OUT(n557),
	.C(n1869),
	.B(n1859),
	.A(n1860));
   INVERTER U1289 (.IN(\mult_19_3/ab[5][4] ),
	.OUT(n1870));
   OAI22 U1290 (.OUT(n1871),
	.D(n1198),
	.C(n1862),
	.B(n561),
	.A(n1872));
   INVERTER U1291 (.IN(\mult_19_3/ab[6][3] ),
	.OUT(n1873));
   OAI21 U1292 (.OUT(n569),
	.C(n1875),
	.B(n1864),
	.A(n1874));
   INVERTER U1293 (.IN(\mult_19_3/ab[5][5] ),
	.OUT(n1876));
   AOI22 U1294 (.A(n557),
	.B(\mult_19_3/ab[4][5] ),
	.C(n1878),
	.D(n1210),
	.OUT(n1877));
   INVERTER U1295 (.IN(\mult_19_3/ab[6][4] ),
	.OUT(n1879));
   OAI21 U1296 (.OUT(n606),
	.C(n1881),
	.B(n1870),
	.A(n1880));
   OAI22 U1297 (.OUT(n608),
	.D(n1213),
	.C(n1873),
	.B(n568),
	.A(n1882));
   NAND2 U1298 (.A(\mult_19_3/ab[0][2] ),
	.B(\mult_19_3/ab[1][1] ),
	.OUT(n1883));
   AOI22 U1299 (.A(\mult_19_3/ab[2][1] ),
	.B(n579),
	.C(n1885),
	.D(n1220),
	.OUT(n1884));
   INVERTER U1300 (.IN(\mult_19_3/ab[3][1] ),
	.OUT(n1886));
   OAI21 U1301 (.OUT(n581),
	.C(n1887),
	.B(n1886),
	.A(n1884));
   OAI22 U1302 (.OUT(n1888),
	.D(n1233),
	.C(n1890),
	.B(n580),
	.A(n1889));
   INVERTER U1303 (.IN(\mult_19_3/ab[5][1] ),
	.OUT(n1891));
   OAI21 U1304 (.OUT(n583),
	.C(n1893),
	.B(n1891),
	.A(n1892));
   OAI22 U1305 (.OUT(n585),
	.D(n1236),
	.C(n1895),
	.B(n582),
	.A(n1894));
   NAND2 U1306 (.A(\mult_19_3/ab[0][1] ),
	.B(\mult_19_3/ab[1][0] ),
	.OUT(n1896));
   AOI22 U1307 (.A(\mult_19_3/ab[2][0] ),
	.B(n587),
	.C(n1898),
	.D(n1229),
	.OUT(n1897));
   INVERTER U1308 (.IN(\mult_19_3/ab[3][0] ),
	.OUT(n1899));
   OAI21 U1309 (.OUT(n589),
	.C(n1900),
	.B(n1899),
	.A(n1897));
   INVERTER U1310 (.IN(\mult_19_3/ab[4][0] ),
	.OUT(n1901));
   OAI22 U1311 (.OUT(n1902),
	.D(n1904),
	.C(n1901),
	.B(n588),
	.A(n1903));
   INVERTER U1312 (.IN(\mult_19_3/ab[5][0] ),
	.OUT(n1905));
   OAI21 U1313 (.OUT(n591),
	.C(n1907),
	.B(n1905),
	.A(n1906));
   INVERTER U1314 (.IN(\mult_19_3/ab[6][0] ),
	.OUT(n1908));
   OAI22 U1315 (.OUT(n593),
	.D(n1910),
	.C(n1908),
	.B(n590),
	.A(n1909));
   INVERTER U1316 (.IN(\mult_19_3/ab[7][7] ),
	.OUT(n99));
   OAI21 U1317 (.OUT(n601),
	.C(n1911),
	.B(n1876),
	.A(n1877));
   AOI22 U1318 (.A(n601),
	.B(\mult_19_3/ab[6][5] ),
	.C(n1912),
	.D(n1239),
	.OUT(n604));
   INVERTER U1319 (.IN(\mult_19_3/ab[7][5] ),
	.OUT(n603));
   OAI22 U1320 (.OUT(n1913),
	.D(n1215),
	.C(n1879),
	.B(n605),
	.A(n1914));
   INVERTER U1321 (.IN(\mult_19_3/ab[7][4] ),
	.OUT(n1915));
   NAND2 U1322 (.A(\mult_19_2/ab[0][3] ),
	.B(\mult_19_2/ab[1][2] ),
	.OUT(n1916));
   AOI22 U1323 (.A(\mult_19_2/ab[2][2] ),
	.B(n628),
	.C(n1918),
	.D(n1260),
	.OUT(n1917));
   NAND2 U1324 (.A(\mult_19_2/ab[1][3] ),
	.B(\mult_19_2/ab[0][4] ),
	.OUT(n622));
   INVERTER U1325 (.IN(\mult_19_2/ab[3][2] ),
	.OUT(n1919));
   OAI21 U1326 (.OUT(n630),
	.C(n1920),
	.B(n1919),
	.A(n1917));
   NAND2 U1327 (.A(\mult_19_2/ab[1][4] ),
	.B(\mult_19_2/ab[0][5] ),
	.OUT(n617));
   INVERTER U1328 (.IN(\mult_19_2/ab[3][3] ),
	.OUT(n1921));
   AOI22 U1329 (.A(n1923),
	.B(\mult_19_2/ab[2][3] ),
	.C(n620),
	.D(n1257),
	.OUT(n1922));
   AOI22 U1330 (.A(n630),
	.B(\mult_19_2/ab[4][2] ),
	.C(n1925),
	.D(n1281),
	.OUT(n1924));
   NAND2 U1331 (.A(\mult_19_2/ab[1][5] ),
	.B(\mult_19_2/ab[0][6] ),
	.OUT(n612));
   INVERTER U1332 (.IN(\mult_19_2/ab[3][4] ),
	.OUT(n1926));
   AOI22 U1333 (.A(n1928),
	.B(\mult_19_2/ab[2][4] ),
	.C(n615),
	.D(n1251),
	.OUT(n1927));
   INVERTER U1334 (.IN(\mult_19_2/ab[4][3] ),
	.OUT(n1929));
   OAI21 U1335 (.OUT(n624),
	.C(n1930),
	.B(n1921),
	.A(n1922));
   INVERTER U1336 (.IN(\mult_19_2/ab[5][2] ),
	.OUT(n1931));
   OAI21 U1337 (.OUT(n632),
	.C(n1932),
	.B(n1931),
	.A(n1924));
   NAND2 U1338 (.A(\mult_19_2/ab[1][6] ),
	.B(\mult_19_2/ab[0][7] ),
	.OUT(n1933));
   INVERTER U1339 (.IN(\mult_19_2/ab[2][6] ),
	.OUT(n1934));
   INVERTER U1340 (.IN(\mult_19_2/ab[1][7] ),
	.OUT(n1935));
   INVERTER U1341 (.IN(\mult_19_2/ab[3][5] ),
	.OUT(n1936));
   AOI22 U1342 (.A(n1938),
	.B(\mult_19_2/ab[2][5] ),
	.C(n610),
	.D(n1250),
	.OUT(n1937));
   INVERTER U1343 (.IN(\mult_19_2/ab[4][4] ),
	.OUT(n1939));
   OAI21 U1344 (.OUT(n619),
	.C(n1940),
	.B(n1926),
	.A(n1927));
   INVERTER U1345 (.IN(\mult_19_2/ab[5][3] ),
	.OUT(n1941));
   OAI22 U1346 (.OUT(n1942),
	.D(n1264),
	.C(n1929),
	.B(n623),
	.A(n1943));
   OAI22 U1347 (.OUT(n634),
	.D(n1284),
	.C(n1945),
	.B(n631),
	.A(n1944));
   OAI21 U1348 (.OUT(n614),
	.C(n1946),
	.B(n1936),
	.A(n1937));
   INVERTER U1349 (.IN(\mult_19_2/ab[5][4] ),
	.OUT(n1947));
   OAI22 U1350 (.OUT(n1948),
	.D(n1255),
	.C(n1939),
	.B(n618),
	.A(n1949));
   INVERTER U1351 (.IN(\mult_19_2/ab[6][3] ),
	.OUT(n1950));
   OAI21 U1352 (.OUT(n626),
	.C(n1952),
	.B(n1941),
	.A(n1951));
   INVERTER U1353 (.IN(\mult_19_2/ab[5][5] ),
	.OUT(n1953));
   AOI22 U1354 (.A(n614),
	.B(\mult_19_2/ab[4][5] ),
	.C(n1955),
	.D(n1267),
	.OUT(n1954));
   INVERTER U1355 (.IN(\mult_19_2/ab[6][4] ),
	.OUT(n1956));
   OAI21 U1356 (.OUT(n663),
	.C(n1958),
	.B(n1947),
	.A(n1957));
   OAI22 U1357 (.OUT(n665),
	.D(n1270),
	.C(n1950),
	.B(n625),
	.A(n1959));
   NAND2 U1358 (.A(\mult_19_2/ab[0][2] ),
	.B(\mult_19_2/ab[1][1] ),
	.OUT(n1960));
   AOI22 U1359 (.A(\mult_19_2/ab[2][1] ),
	.B(n636),
	.C(n1962),
	.D(n1277),
	.OUT(n1961));
   INVERTER U1360 (.IN(\mult_19_2/ab[3][1] ),
	.OUT(n1963));
   OAI21 U1361 (.OUT(n638),
	.C(n1964),
	.B(n1963),
	.A(n1961));
   OAI22 U1362 (.OUT(n1965),
	.D(n1290),
	.C(n1967),
	.B(n637),
	.A(n1966));
   INVERTER U1363 (.IN(\mult_19_2/ab[5][1] ),
	.OUT(n1968));
   OAI21 U1364 (.OUT(n640),
	.C(n1970),
	.B(n1968),
	.A(n1969));
   OAI22 U1365 (.OUT(n642),
	.D(n1293),
	.C(n1972),
	.B(n639),
	.A(n1971));
   NAND2 U1366 (.A(\mult_19_2/ab[0][1] ),
	.B(\mult_19_2/ab[1][0] ),
	.OUT(n1973));
   AOI22 U1367 (.A(\mult_19_2/ab[2][0] ),
	.B(n644),
	.C(n1975),
	.D(n1286),
	.OUT(n1974));
   INVERTER U1368 (.IN(\mult_19_2/ab[3][0] ),
	.OUT(n1976));
   OAI21 U1369 (.OUT(n646),
	.C(n1977),
	.B(n1976),
	.A(n1974));
   INVERTER U1370 (.IN(\mult_19_2/ab[4][0] ),
	.OUT(n1978));
   OAI22 U1371 (.OUT(n1979),
	.D(n1981),
	.C(n1978),
	.B(n645),
	.A(n1980));
   INVERTER U1372 (.IN(\mult_19_2/ab[5][0] ),
	.OUT(n1982));
   OAI21 U1373 (.OUT(n648),
	.C(n1984),
	.B(n1982),
	.A(n1983));
   INVERTER U1374 (.IN(\mult_19_2/ab[6][0] ),
	.OUT(n1985));
   OAI22 U1375 (.OUT(n650),
	.D(n1987),
	.C(n1985),
	.B(n647),
	.A(n1986));
   INVERTER U1376 (.IN(\mult_19_2/ab[7][7] ),
	.OUT(n83));
   OAI21 U1377 (.OUT(n658),
	.C(n1988),
	.B(n1953),
	.A(n1954));
   AOI22 U1378 (.A(n658),
	.B(\mult_19_2/ab[6][5] ),
	.C(n1989),
	.D(n1296),
	.OUT(n661));
   INVERTER U1379 (.IN(\mult_19_2/ab[7][5] ),
	.OUT(n660));
   OAI22 U1380 (.OUT(n1990),
	.D(n1272),
	.C(n1956),
	.B(n662),
	.A(n1991));
   INVERTER U1381 (.IN(\mult_19_2/ab[7][4] ),
	.OUT(n1992));
   NAND2 U1382 (.A(\mult_19/ab[0][3] ),
	.B(\mult_19/ab[1][2] ),
	.OUT(n1993));
   AOI22 U1383 (.A(\mult_19/ab[2][2] ),
	.B(n685),
	.C(n1995),
	.D(n1317),
	.OUT(n1994));
   NAND2 U1384 (.A(\mult_19/ab[1][3] ),
	.B(\mult_19/ab[0][4] ),
	.OUT(n679));
   INVERTER U1385 (.IN(\mult_19/ab[3][2] ),
	.OUT(n1996));
   OAI21 U1386 (.OUT(n687),
	.C(n1997),
	.B(n1996),
	.A(n1994));
   NAND2 U1387 (.A(\mult_19/ab[1][4] ),
	.B(\mult_19/ab[0][5] ),
	.OUT(n674));
   INVERTER U1388 (.IN(\mult_19/ab[3][3] ),
	.OUT(n1998));
   AOI22 U1389 (.A(n2000),
	.B(\mult_19/ab[2][3] ),
	.C(n677),
	.D(n1314),
	.OUT(n1999));
   AOI22 U1390 (.A(n687),
	.B(\mult_19/ab[4][2] ),
	.C(n2002),
	.D(n1338),
	.OUT(n2001));
   NAND2 U1391 (.A(\mult_19/ab[1][5] ),
	.B(\mult_19/ab[0][6] ),
	.OUT(n669));
   INVERTER U1392 (.IN(\mult_19/ab[3][4] ),
	.OUT(n2003));
   AOI22 U1393 (.A(n2005),
	.B(\mult_19/ab[2][4] ),
	.C(n672),
	.D(n1308),
	.OUT(n2004));
   INVERTER U1394 (.IN(\mult_19/ab[4][3] ),
	.OUT(n2006));
   OAI21 U1395 (.OUT(n681),
	.C(n2007),
	.B(n1998),
	.A(n1999));
   INVERTER U1396 (.IN(\mult_19/ab[5][2] ),
	.OUT(n2008));
   OAI21 U1397 (.OUT(n689),
	.C(n2009),
	.B(n2008),
	.A(n2001));
   NAND2 U1398 (.A(\mult_19/ab[1][6] ),
	.B(\mult_19/ab[0][7] ),
	.OUT(n2010));
   INVERTER U1399 (.IN(\mult_19/ab[2][6] ),
	.OUT(n2011));
   INVERTER U1400 (.IN(\mult_19/ab[1][7] ),
	.OUT(n2012));
   INVERTER U1401 (.IN(\mult_19/ab[3][5] ),
	.OUT(n2013));
   AOI22 U1402 (.A(n2015),
	.B(\mult_19/ab[2][5] ),
	.C(n667),
	.D(n1307),
	.OUT(n2014));
   INVERTER U1403 (.IN(\mult_19/ab[4][4] ),
	.OUT(n2016));
   OAI21 U1404 (.OUT(n676),
	.C(n2017),
	.B(n2003),
	.A(n2004));
   INVERTER U1405 (.IN(\mult_19/ab[5][3] ),
	.OUT(n2018));
   OAI22 U1406 (.OUT(n2019),
	.D(n1321),
	.C(n2006),
	.B(n680),
	.A(n2020));
   OAI22 U1407 (.OUT(n691),
	.D(n1341),
	.C(n2022),
	.B(n688),
	.A(n2021));
   OAI21 U1408 (.OUT(n671),
	.C(n2023),
	.B(n2013),
	.A(n2014));
   INVERTER U1409 (.IN(\mult_19/ab[5][4] ),
	.OUT(n2024));
   OAI22 U1410 (.OUT(n2025),
	.D(n1312),
	.C(n2016),
	.B(n675),
	.A(n2026));
   INVERTER U1411 (.IN(\mult_19/ab[6][3] ),
	.OUT(n2027));
   OAI21 U1412 (.OUT(n683),
	.C(n2029),
	.B(n2018),
	.A(n2028));
   INVERTER U1413 (.IN(\mult_19/ab[5][5] ),
	.OUT(n2030));
   AOI22 U1414 (.A(n671),
	.B(\mult_19/ab[4][5] ),
	.C(n2032),
	.D(n1324),
	.OUT(n2031));
   INVERTER U1415 (.IN(\mult_19/ab[6][4] ),
	.OUT(n2033));
   OAI21 U1416 (.OUT(n720),
	.C(n2035),
	.B(n2024),
	.A(n2034));
   OAI22 U1417 (.OUT(n722),
	.D(n1327),
	.C(n2027),
	.B(n682),
	.A(n2036));
   NAND2 U1418 (.A(\mult_19/ab[0][2] ),
	.B(\mult_19/ab[1][1] ),
	.OUT(n2037));
   AOI22 U1419 (.A(\mult_19/ab[2][1] ),
	.B(n693),
	.C(n2039),
	.D(n1334),
	.OUT(n2038));
   INVERTER U1420 (.IN(\mult_19/ab[3][1] ),
	.OUT(n2040));
   OAI21 U1421 (.OUT(n695),
	.C(n2041),
	.B(n2040),
	.A(n2038));
   OAI22 U1422 (.OUT(n2042),
	.D(n1347),
	.C(n2044),
	.B(n694),
	.A(n2043));
   INVERTER U1423 (.IN(\mult_19/ab[5][1] ),
	.OUT(n2045));
   OAI21 U1424 (.OUT(n697),
	.C(n2047),
	.B(n2045),
	.A(n2046));
   OAI22 U1425 (.OUT(n699),
	.D(n1350),
	.C(n2049),
	.B(n696),
	.A(n2048));
   NAND2 U1426 (.A(\mult_19/ab[0][1] ),
	.B(\mult_19/ab[1][0] ),
	.OUT(n2050));
   AOI22 U1427 (.A(\mult_19/ab[2][0] ),
	.B(n701),
	.C(n2052),
	.D(n1343),
	.OUT(n2051));
   INVERTER U1428 (.IN(\mult_19/ab[3][0] ),
	.OUT(n2053));
   OAI21 U1429 (.OUT(n703),
	.C(n2054),
	.B(n2053),
	.A(n2051));
   INVERTER U1430 (.IN(\mult_19/ab[4][0] ),
	.OUT(n2055));
   OAI22 U1431 (.OUT(n2056),
	.D(n2058),
	.C(n2055),
	.B(n702),
	.A(n2057));
   INVERTER U1432 (.IN(\mult_19/ab[5][0] ),
	.OUT(n2059));
   OAI21 U1433 (.OUT(n705),
	.C(n2061),
	.B(n2059),
	.A(n2060));
   INVERTER U1434 (.IN(\mult_19/ab[6][0] ),
	.OUT(n2062));
   OAI22 U1435 (.OUT(n707),
	.D(n2064),
	.C(n2062),
	.B(n704),
	.A(n2063));
   INVERTER U1436 (.IN(\mult_19/ab[7][7] ),
	.OUT(n67));
   OAI21 U1437 (.OUT(n715),
	.C(n2065),
	.B(n2030),
	.A(n2031));
   AOI22 U1438 (.A(n715),
	.B(\mult_19/ab[6][5] ),
	.C(n2066),
	.D(n1353),
	.OUT(n718));
   INVERTER U1439 (.IN(\mult_19/ab[7][5] ),
	.OUT(n717));
   OAI22 U1440 (.OUT(n2067),
	.D(n1329),
	.C(n2033),
	.B(n719),
	.A(n2068));
   INVERTER U1441 (.IN(\mult_19/ab[7][4] ),
	.OUT(n2069));
   NAND2 U1442 (.A(N1),
	.B(N17),
	.OUT(n2070));
   INVERTER U1443 (.IN(N31),
	.OUT(n2071));
   INVERTER U1444 (.IN(N15),
	.OUT(n2072));
   NAND2 U1445 (.A(N49),
	.B(n1364),
	.OUT(n2073));
   AOI22 U1446 (.A(n737),
	.B(n736),
	.C(n2074),
	.D(n1365),
	.OUT(n740));
   AOI22 U1447 (.A(n2076),
	.B(N51),
	.C(n738),
	.D(n2077),
	.OUT(n2075));
   INVERTER U1448 (.IN(N52),
	.OUT(n2078));
   OAI21 U1449 (.OUT(n742),
	.C(n2079),
	.B(n2078),
	.A(n2075));
   AOI22 U1450 (.A(n742),
	.B(N53),
	.C(n2080),
	.D(n2081),
	.OUT(n745));
   INVERTER U1451 (.IN(N54),
	.OUT(n744));
   OAI22 U1452 (.OUT(n2082),
	.D(n2084),
	.C(n744),
	.B(n2083),
	.A(n745));
   INVERTER U1453 (.IN(N55),
	.OUT(n2085));
   OAI21 U1454 (.OUT(n747),
	.C(n2087),
	.B(n2085),
	.A(n2086));
   INVERTER U1455 (.IN(N56),
	.OUT(n2088));
   OAI22 U1456 (.OUT(n749),
	.D(n2090),
	.C(n2088),
	.B(n746),
	.A(n2089));
   AOI22 U1457 (.A(n749),
	.B(N57),
	.C(n2091),
	.D(n2092),
	.OUT(n752));
   INVERTER U1458 (.IN(N58),
	.OUT(n751));
   OAI22 U1459 (.OUT(n754),
	.D(n2094),
	.C(n751),
	.B(n2093),
	.A(n752));
   AOI22 U1460 (.A(n754),
	.B(N59),
	.C(n2095),
	.D(n2096),
	.OUT(n757));
   INVERTER U1461 (.IN(N60),
	.OUT(n756));
   OAI22 U1462 (.OUT(n759),
	.D(n2098),
	.C(n756),
	.B(n2097),
	.A(n757));
   AOI22 U1463 (.A(n759),
	.B(N61),
	.C(n2099),
	.D(n2100),
	.OUT(n762));
   INVERTER U1464 (.IN(N62),
	.OUT(n761));
   OAI22 U1465 (.OUT(n764),
	.D(n2102),
	.C(n761),
	.B(n2101),
	.A(n762));
   INVERTER U1466 (.IN(N63),
	.OUT(n2103));
   NAND2 U1467 (.A(N161),
	.B(N177),
	.OUT(n2104));
   INVERTER U1468 (.IN(N191),
	.OUT(n2105));
   INVERTER U1469 (.IN(N175),
	.OUT(n2106));
   NAND2 U1470 (.A(N209),
	.B(n1369),
	.OUT(n2107));
   AOI22 U1471 (.A(n779),
	.B(n778),
	.C(n2108),
	.D(n1370),
	.OUT(n782));
   AOI22 U1472 (.A(n2110),
	.B(N211),
	.C(n780),
	.D(n2111),
	.OUT(n2109));
   INVERTER U1473 (.IN(N212),
	.OUT(n2112));
   OAI21 U1474 (.OUT(n784),
	.C(n2113),
	.B(n2112),
	.A(n2109));
   AOI22 U1475 (.A(n784),
	.B(N213),
	.C(n2114),
	.D(n2115),
	.OUT(n787));
   INVERTER U1476 (.IN(N214),
	.OUT(n786));
   OAI22 U1477 (.OUT(n2116),
	.D(n2118),
	.C(n786),
	.B(n2117),
	.A(n787));
   INVERTER U1478 (.IN(N215),
	.OUT(n2119));
   OAI21 U1479 (.OUT(n789),
	.C(n2121),
	.B(n2119),
	.A(n2120));
   INVERTER U1480 (.IN(N216),
	.OUT(n2122));
   OAI22 U1481 (.OUT(n791),
	.D(n2124),
	.C(n2122),
	.B(n788),
	.A(n2123));
   AOI22 U1482 (.A(n791),
	.B(N217),
	.C(n2125),
	.D(n2126),
	.OUT(n794));
   INVERTER U1483 (.IN(N218),
	.OUT(n793));
   OAI22 U1484 (.OUT(n796),
	.D(n2128),
	.C(n793),
	.B(n2127),
	.A(n794));
   AOI22 U1485 (.A(n796),
	.B(N219),
	.C(n2129),
	.D(n2130),
	.OUT(n799));
   INVERTER U1486 (.IN(N220),
	.OUT(n798));
   OAI22 U1487 (.OUT(n801),
	.D(n2132),
	.C(n798),
	.B(n2131),
	.A(n799));
   AOI22 U1488 (.A(n801),
	.B(N221),
	.C(n2133),
	.D(n2134),
	.OUT(n804));
   INVERTER U1489 (.IN(N222),
	.OUT(n803));
   OAI22 U1490 (.OUT(n806),
	.D(n2136),
	.C(n803),
	.B(n2135),
	.A(n804));
   INVERTER U1491 (.IN(N223),
	.OUT(n2137));
   NAND2 U1492 (.A(N81),
	.B(N97),
	.OUT(n2138));
   INVERTER U1493 (.IN(N111),
	.OUT(n2139));
   INVERTER U1494 (.IN(N95),
	.OUT(n2140));
   NAND2 U1495 (.A(N129),
	.B(n1374),
	.OUT(n2141));
   AOI22 U1496 (.A(n821),
	.B(n820),
	.C(n2142),
	.D(n1375),
	.OUT(n824));
   AOI22 U1497 (.A(n2144),
	.B(N131),
	.C(n822),
	.D(n2145),
	.OUT(n2143));
   INVERTER U1498 (.IN(N132),
	.OUT(n2146));
   OAI21 U1499 (.OUT(n826),
	.C(n2147),
	.B(n2146),
	.A(n2143));
   AOI22 U1500 (.A(n826),
	.B(N133),
	.C(n2148),
	.D(n2149),
	.OUT(n829));
   INVERTER U1501 (.IN(N134),
	.OUT(n828));
   OAI22 U1502 (.OUT(n2150),
	.D(n2152),
	.C(n828),
	.B(n2151),
	.A(n829));
   INVERTER U1503 (.IN(N135),
	.OUT(n2153));
   OAI21 U1504 (.OUT(n831),
	.C(n2155),
	.B(n2153),
	.A(n2154));
   INVERTER U1505 (.IN(N136),
	.OUT(n2156));
   OAI22 U1506 (.OUT(n833),
	.D(n2158),
	.C(n2156),
	.B(n830),
	.A(n2157));
   AOI22 U1507 (.A(n833),
	.B(N137),
	.C(n2159),
	.D(n2160),
	.OUT(n836));
   INVERTER U1508 (.IN(N138),
	.OUT(n835));
   OAI22 U1509 (.OUT(n838),
	.D(n2162),
	.C(n835),
	.B(n2161),
	.A(n836));
   AOI22 U1510 (.A(n838),
	.B(N139),
	.C(n2163),
	.D(n2164),
	.OUT(n841));
   INVERTER U1511 (.IN(N140),
	.OUT(n840));
   OAI22 U1512 (.OUT(n843),
	.D(n2166),
	.C(n840),
	.B(n2165),
	.A(n841));
   AOI22 U1513 (.A(n843),
	.B(N141),
	.C(n2167),
	.D(n2168),
	.OUT(n846));
   INVERTER U1514 (.IN(N142),
	.OUT(n845));
   OAI22 U1515 (.OUT(n848),
	.D(n2170),
	.C(n845),
	.B(n2169),
	.A(n846));
   INVERTER U1516 (.IN(N143),
	.OUT(n2171));
   XOR2 U1517 (.A(n202),
	.B(n203),
	.OUT(\mult_21_3/A1[9] ));
   XOR2 U1518 (.A(n206),
	.B(n207),
	.OUT(\mult_21_3/A1[7] ));
   XOR2 U1519 (.A(n208),
	.B(n209),
	.OUT(\mult_21_3/A1[6] ));
   XOR2 U1520 (.A(n1448),
	.B(n2172),
	.OUT(\mult_21_3/A1[4] ));
   XOR2 U1521 (.A(n1442),
	.B(n2173),
	.OUT(\mult_21_3/A1[2] ));
   XOR2 U1522 (.A(n197),
	.B(n198),
	.OUT(\mult_21_3/A1[11] ));
   XOR2 U1523 (.A(n887),
	.B(n2174),
	.OUT(\mult_21_3/A1[0] ));
   XOR2 U1524 (.A(n186),
	.B(n187),
	.OUT(\mult_21_2/A1[9] ));
   XOR2 U1525 (.A(n190),
	.B(n191),
	.OUT(\mult_21_2/A1[7] ));
   XOR2 U1526 (.A(n192),
	.B(n193),
	.OUT(\mult_21_2/A1[6] ));
   XOR2 U1527 (.A(n1525),
	.B(n2175),
	.OUT(\mult_21_2/A1[4] ));
   XOR2 U1528 (.A(n1519),
	.B(n2176),
	.OUT(\mult_21_2/A1[2] ));
   XOR2 U1529 (.A(n181),
	.B(n182),
	.OUT(\mult_21_2/A1[11] ));
   XOR2 U1530 (.A(n944),
	.B(n2177),
	.OUT(\mult_21_2/A1[0] ));
   XOR2 U1531 (.A(n170),
	.B(n171),
	.OUT(\mult_21/A1[9] ));
   XOR2 U1532 (.A(n174),
	.B(n175),
	.OUT(\mult_21/A1[7] ));
   XOR2 U1533 (.A(n176),
	.B(n177),
	.OUT(\mult_21/A1[6] ));
   XOR2 U1534 (.A(n1602),
	.B(n2178),
	.OUT(\mult_21/A1[4] ));
   XOR2 U1535 (.A(n1596),
	.B(n2179),
	.OUT(\mult_21/A1[2] ));
   XOR2 U1536 (.A(n165),
	.B(n166),
	.OUT(\mult_21/A1[11] ));
   XOR2 U1537 (.A(n1001),
	.B(n2180),
	.OUT(\mult_21/A1[0] ));
   XOR2 U1538 (.A(n154),
	.B(n155),
	.OUT(\mult_20_3/A1[9] ));
   XOR2 U1539 (.A(n158),
	.B(n159),
	.OUT(\mult_20_3/A1[7] ));
   XOR2 U1540 (.A(n160),
	.B(n161),
	.OUT(\mult_20_3/A1[6] ));
   XOR2 U1541 (.A(n1679),
	.B(n2181),
	.OUT(\mult_20_3/A1[4] ));
   XOR2 U1542 (.A(n1673),
	.B(n2182),
	.OUT(\mult_20_3/A1[2] ));
   XOR2 U1543 (.A(n149),
	.B(n150),
	.OUT(\mult_20_3/A1[11] ));
   XOR2 U1544 (.A(n1058),
	.B(n2183),
	.OUT(\mult_20_3/A1[0] ));
   XOR2 U1545 (.A(n138),
	.B(n139),
	.OUT(\mult_20_2/A1[9] ));
   XOR2 U1546 (.A(n142),
	.B(n143),
	.OUT(\mult_20_2/A1[7] ));
   XOR2 U1547 (.A(n144),
	.B(n145),
	.OUT(\mult_20_2/A1[6] ));
   XOR2 U1548 (.A(n1756),
	.B(n2184),
	.OUT(\mult_20_2/A1[4] ));
   XOR2 U1549 (.A(n1750),
	.B(n2185),
	.OUT(\mult_20_2/A1[2] ));
   XOR2 U1550 (.A(n133),
	.B(n134),
	.OUT(\mult_20_2/A1[11] ));
   XOR2 U1551 (.A(n1115),
	.B(n2186),
	.OUT(\mult_20_2/A1[0] ));
   XOR2 U1552 (.A(n122),
	.B(n123),
	.OUT(\mult_20/A1[9] ));
   XOR2 U1553 (.A(n126),
	.B(n127),
	.OUT(\mult_20/A1[7] ));
   XOR2 U1554 (.A(n128),
	.B(n129),
	.OUT(\mult_20/A1[6] ));
   XOR2 U1555 (.A(n1833),
	.B(n2187),
	.OUT(\mult_20/A1[4] ));
   XOR2 U1556 (.A(n1827),
	.B(n2188),
	.OUT(\mult_20/A1[2] ));
   XOR2 U1557 (.A(n117),
	.B(n118),
	.OUT(\mult_20/A1[11] ));
   XOR2 U1558 (.A(n1172),
	.B(n2189),
	.OUT(\mult_20/A1[0] ));
   XOR2 U1559 (.A(n106),
	.B(n107),
	.OUT(\mult_19_3/A1[9] ));
   XOR2 U1560 (.A(n110),
	.B(n111),
	.OUT(\mult_19_3/A1[7] ));
   XOR2 U1561 (.A(n112),
	.B(n113),
	.OUT(\mult_19_3/A1[6] ));
   XOR2 U1562 (.A(n1910),
	.B(n2190),
	.OUT(\mult_19_3/A1[4] ));
   XOR2 U1563 (.A(n1904),
	.B(n2191),
	.OUT(\mult_19_3/A1[2] ));
   XOR2 U1564 (.A(n101),
	.B(n102),
	.OUT(\mult_19_3/A1[11] ));
   XOR2 U1565 (.A(n1229),
	.B(n2192),
	.OUT(\mult_19_3/A1[0] ));
   XOR2 U1566 (.A(n90),
	.B(n91),
	.OUT(\mult_19_2/A1[9] ));
   XOR2 U1567 (.A(n94),
	.B(n95),
	.OUT(\mult_19_2/A1[7] ));
   XOR2 U1568 (.A(n96),
	.B(n97),
	.OUT(\mult_19_2/A1[6] ));
   XOR2 U1569 (.A(n1987),
	.B(n2193),
	.OUT(\mult_19_2/A1[4] ));
   XOR2 U1570 (.A(n1981),
	.B(n2194),
	.OUT(\mult_19_2/A1[2] ));
   XOR2 U1571 (.A(n85),
	.B(n86),
	.OUT(\mult_19_2/A1[11] ));
   XOR2 U1572 (.A(n1286),
	.B(n2195),
	.OUT(\mult_19_2/A1[0] ));
   XOR2 U1573 (.A(n74),
	.B(n75),
	.OUT(\mult_19/A1[9] ));
   XOR2 U1574 (.A(n78),
	.B(n79),
	.OUT(\mult_19/A1[7] ));
   XOR2 U1575 (.A(n80),
	.B(n81),
	.OUT(\mult_19/A1[6] ));
   XOR2 U1576 (.A(n2064),
	.B(n2196),
	.OUT(\mult_19/A1[4] ));
   XOR2 U1577 (.A(n2058),
	.B(n2197),
	.OUT(\mult_19/A1[2] ));
   XOR2 U1578 (.A(n69),
	.B(n70),
	.OUT(\mult_19/A1[11] ));
   XOR2 U1579 (.A(n1343),
	.B(n2198),
	.OUT(\mult_19/A1[0] ));
   XOR2 U1580 (.A(n2199),
	.B(n2200),
	.OUT(N80));
   XOR2 U1581 (.A(n2201),
	.B(n2202),
	.OUT(N79));
   XOR2 U1582 (.A(n2102),
	.B(n2203),
	.OUT(N78));
   XOR2 U1583 (.A(n2100),
	.B(n2204),
	.OUT(N77));
   XOR2 U1584 (.A(n2098),
	.B(n2205),
	.OUT(N76));
   XOR2 U1585 (.A(n2096),
	.B(n2206),
	.OUT(N75));
   XOR2 U1586 (.A(n2094),
	.B(n2207),
	.OUT(N74));
   XOR2 U1587 (.A(n2092),
	.B(n2208),
	.OUT(N73));
   XOR2 U1588 (.A(n2090),
	.B(n2209),
	.OUT(N72));
   XOR2 U1589 (.A(n2210),
	.B(n2211),
	.OUT(N71));
   XOR2 U1590 (.A(n2084),
	.B(n2212),
	.OUT(N70));
   XOR2 U1591 (.A(n2081),
	.B(n2213),
	.OUT(N69));
   XOR2 U1592 (.A(n2214),
	.B(n2215),
	.OUT(N68));
   XOR2 U1593 (.A(n2216),
	.B(n2217),
	.OUT(N67));
   XOR2 U1594 (.A(n1365),
	.B(n2218),
	.OUT(N66));
   XOR2 U1595 (.A(N49),
	.B(n1364),
	.OUT(N65));
   XOR2 U1596 (.A(n2219),
	.B(n2220),
	.OUT(N240));
   XOR2 U1597 (.A(n2221),
	.B(n2222),
	.OUT(N239));
   XOR2 U1598 (.A(n2136),
	.B(n2223),
	.OUT(N238));
   XOR2 U1599 (.A(n2134),
	.B(n2224),
	.OUT(N237));
   XOR2 U1600 (.A(n2132),
	.B(n2225),
	.OUT(N236));
   XOR2 U1601 (.A(n2130),
	.B(n2226),
	.OUT(N235));
   XOR2 U1602 (.A(n2128),
	.B(n2227),
	.OUT(N234));
   XOR2 U1603 (.A(n2126),
	.B(n2228),
	.OUT(N233));
   XOR2 U1604 (.A(n2124),
	.B(n2229),
	.OUT(N232));
   XOR2 U1605 (.A(n2230),
	.B(n2231),
	.OUT(N231));
   XOR2 U1606 (.A(n2118),
	.B(n2232),
	.OUT(N230));
   XOR2 U1607 (.A(n2115),
	.B(n2233),
	.OUT(N229));
   XOR2 U1608 (.A(n2234),
	.B(n2235),
	.OUT(N228));
   XOR2 U1609 (.A(n2236),
	.B(n2237),
	.OUT(N227));
   XOR2 U1610 (.A(n1370),
	.B(n2238),
	.OUT(N226));
   XOR2 U1611 (.A(N209),
	.B(n1369),
	.OUT(N225));
   XOR2 U1612 (.A(n2239),
	.B(n2240),
	.OUT(N160));
   XOR2 U1613 (.A(n2241),
	.B(n2242),
	.OUT(N159));
   XOR2 U1614 (.A(n2170),
	.B(n2243),
	.OUT(N158));
   XOR2 U1615 (.A(n2168),
	.B(n2244),
	.OUT(N157));
   XOR2 U1616 (.A(n2166),
	.B(n2245),
	.OUT(N156));
   XOR2 U1617 (.A(n2164),
	.B(n2246),
	.OUT(N155));
   XOR2 U1618 (.A(n2162),
	.B(n2247),
	.OUT(N154));
   XOR2 U1619 (.A(n2160),
	.B(n2248),
	.OUT(N153));
   XOR2 U1620 (.A(n2158),
	.B(n2249),
	.OUT(N152));
   XOR2 U1621 (.A(n2250),
	.B(n2251),
	.OUT(N151));
   XOR2 U1622 (.A(n2152),
	.B(n2252),
	.OUT(N150));
   XOR2 U1623 (.A(n2149),
	.B(n2253),
	.OUT(N149));
   XOR2 U1624 (.A(n2254),
	.B(n2255),
	.OUT(N148));
   XOR2 U1625 (.A(n2256),
	.B(n2257),
	.OUT(N147));
   XOR2 U1626 (.A(n1375),
	.B(n2258),
	.OUT(N146));
   XOR2 U1627 (.A(N129),
	.B(n1374),
	.OUT(N145));
   XOR2 U1628 (.A(n1384),
	.B(\mult_21_3/ab[2][3] ),
	.OUT(n863));
   XOR2 U1629 (.A(n1389),
	.B(\mult_21_3/ab[2][4] ),
	.OUT(n860));
   XOR2 U1630 (.A(n1382),
	.B(n2260),
	.OUT(n2259));
   XOR2 U1631 (.A(n1399),
	.B(\mult_21_3/ab[2][5] ),
	.OUT(n854));
   XOR2 U1632 (.A(n1387),
	.B(n2262),
	.OUT(n2261));
   XOR2 U1633 (.A(n1390),
	.B(n225),
	.OUT(n866));
   XOR2 U1634 (.A(n1394),
	.B(n1395),
	.OUT(n850));
   XOR2 U1635 (.A(n1397),
	.B(n2264),
	.OUT(n2263));
   XOR2 U1636 (.A(n1400),
	.B(n220),
	.OUT(n857));
   XOR2 U1637 (.A(n1402),
	.B(n1403),
	.OUT(n2265));
   XOR2 U1638 (.A(\mult_21_3/ab[4][5] ),
	.B(n215),
	.OUT(n869));
   XOR2 U1639 (.A(n1408),
	.B(n1409),
	.OUT(n2266));
   XOR2 U1640 (.A(n1411),
	.B(n227),
	.OUT(n872));
   XOR2 U1641 (.A(n1414),
	.B(n2267),
	.OUT(n875));
   XOR2 U1642 (.A(n1417),
	.B(n264),
	.OUT(n2268));
   XOR2 U1643 (.A(\mult_21_3/ab[7][3] ),
	.B(n266),
	.OUT(n877));
   XOR2 U1644 (.A(n229),
	.B(\mult_21_3/ab[2][2] ),
	.OUT(n880));
   XOR2 U1645 (.A(n1380),
	.B(n2270),
	.OUT(n2269));
   XOR2 U1646 (.A(\mult_21_3/ab[4][2] ),
	.B(n231),
	.OUT(n883));
   XOR2 U1647 (.A(n1392),
	.B(n2272),
	.OUT(n2271));
   XOR2 U1648 (.A(\mult_21_3/ab[6][2] ),
	.B(n233),
	.OUT(n886));
   XOR2 U1649 (.A(\mult_21_3/ab[7][2] ),
	.B(n235),
	.OUT(n2273));
   XOR2 U1650 (.A(n237),
	.B(\mult_21_3/ab[2][1] ),
	.OUT(n889));
   XOR2 U1651 (.A(n1424),
	.B(n2275),
	.OUT(n2274));
   XOR2 U1652 (.A(\mult_21_3/ab[4][1] ),
	.B(n239),
	.OUT(n892));
   XOR2 U1653 (.A(n1429),
	.B(n1426),
	.OUT(n2276));
   XOR2 U1654 (.A(\mult_21_3/ab[6][1] ),
	.B(n241),
	.OUT(n895));
   XOR2 U1655 (.A(\mult_21_3/ab[7][1] ),
	.B(n243),
	.OUT(n2277));
   XOR2 U1656 (.A(\mult_21_3/ab[6][5] ),
	.B(n259),
	.OUT(n898));
   XOR2 U1657 (.A(\mult_21_3/ab[7][5] ),
	.B(n262),
	.OUT(n900));
   XOR2 U1658 (.A(\mult_21_3/ab[7][4] ),
	.B(n2279),
	.OUT(n2278));
   XOR2 U1659 (.A(\mult_21_3/ab[7][0] ),
	.B(n251),
	.OUT(n902));
   XOR2 U1660 (.A(n1446),
	.B(n249),
	.OUT(n2172));
   XOR2 U1661 (.A(n1443),
	.B(n1440),
	.OUT(n903));
   XOR2 U1662 (.A(n1439),
	.B(n247),
	.OUT(n2173));
   XOR2 U1663 (.A(n1437),
	.B(n2280),
	.OUT(n905));
   XOR2 U1664 (.A(n245),
	.B(\mult_21_3/ab[2][0] ),
	.OUT(n2174));
   XOR2 U1665 (.A(n1461),
	.B(\mult_21_2/ab[2][3] ),
	.OUT(n920));
   XOR2 U1666 (.A(n1466),
	.B(\mult_21_2/ab[2][4] ),
	.OUT(n917));
   XOR2 U1667 (.A(n1459),
	.B(n2282),
	.OUT(n2281));
   XOR2 U1668 (.A(n1476),
	.B(\mult_21_2/ab[2][5] ),
	.OUT(n911));
   XOR2 U1669 (.A(n1464),
	.B(n2284),
	.OUT(n2283));
   XOR2 U1670 (.A(n1467),
	.B(n282),
	.OUT(n923));
   XOR2 U1671 (.A(n1471),
	.B(n1472),
	.OUT(n907));
   XOR2 U1672 (.A(n1474),
	.B(n2286),
	.OUT(n2285));
   XOR2 U1673 (.A(n1477),
	.B(n277),
	.OUT(n914));
   XOR2 U1674 (.A(n1479),
	.B(n1480),
	.OUT(n2287));
   XOR2 U1675 (.A(\mult_21_2/ab[4][5] ),
	.B(n272),
	.OUT(n926));
   XOR2 U1676 (.A(n1485),
	.B(n1486),
	.OUT(n2288));
   XOR2 U1677 (.A(n1488),
	.B(n284),
	.OUT(n929));
   XOR2 U1678 (.A(n1491),
	.B(n2289),
	.OUT(n932));
   XOR2 U1679 (.A(n1494),
	.B(n321),
	.OUT(n2290));
   XOR2 U1680 (.A(\mult_21_2/ab[7][3] ),
	.B(n323),
	.OUT(n934));
   XOR2 U1681 (.A(n286),
	.B(\mult_21_2/ab[2][2] ),
	.OUT(n937));
   XOR2 U1682 (.A(n1457),
	.B(n2292),
	.OUT(n2291));
   XOR2 U1683 (.A(\mult_21_2/ab[4][2] ),
	.B(n288),
	.OUT(n940));
   XOR2 U1684 (.A(n1469),
	.B(n2294),
	.OUT(n2293));
   XOR2 U1685 (.A(\mult_21_2/ab[6][2] ),
	.B(n290),
	.OUT(n943));
   XOR2 U1686 (.A(\mult_21_2/ab[7][2] ),
	.B(n292),
	.OUT(n2295));
   XOR2 U1687 (.A(n294),
	.B(\mult_21_2/ab[2][1] ),
	.OUT(n946));
   XOR2 U1688 (.A(n1501),
	.B(n2297),
	.OUT(n2296));
   XOR2 U1689 (.A(\mult_21_2/ab[4][1] ),
	.B(n296),
	.OUT(n949));
   XOR2 U1690 (.A(n1506),
	.B(n1503),
	.OUT(n2298));
   XOR2 U1691 (.A(\mult_21_2/ab[6][1] ),
	.B(n298),
	.OUT(n952));
   XOR2 U1692 (.A(\mult_21_2/ab[7][1] ),
	.B(n300),
	.OUT(n2299));
   XOR2 U1693 (.A(\mult_21_2/ab[6][5] ),
	.B(n316),
	.OUT(n955));
   XOR2 U1694 (.A(\mult_21_2/ab[7][5] ),
	.B(n319),
	.OUT(n957));
   XOR2 U1695 (.A(\mult_21_2/ab[7][4] ),
	.B(n2301),
	.OUT(n2300));
   XOR2 U1696 (.A(\mult_21_2/ab[7][0] ),
	.B(n308),
	.OUT(n959));
   XOR2 U1697 (.A(n1523),
	.B(n306),
	.OUT(n2175));
   XOR2 U1698 (.A(n1520),
	.B(n1517),
	.OUT(n960));
   XOR2 U1699 (.A(n1516),
	.B(n304),
	.OUT(n2176));
   XOR2 U1700 (.A(n1514),
	.B(n2302),
	.OUT(n962));
   XOR2 U1701 (.A(n302),
	.B(\mult_21_2/ab[2][0] ),
	.OUT(n2177));
   XOR2 U1702 (.A(n1538),
	.B(\mult_21/ab[2][3] ),
	.OUT(n977));
   XOR2 U1703 (.A(n1543),
	.B(\mult_21/ab[2][4] ),
	.OUT(n974));
   XOR2 U1704 (.A(n1536),
	.B(n2304),
	.OUT(n2303));
   XOR2 U1705 (.A(n1553),
	.B(\mult_21/ab[2][5] ),
	.OUT(n968));
   XOR2 U1706 (.A(n1541),
	.B(n2306),
	.OUT(n2305));
   XOR2 U1707 (.A(n1544),
	.B(n339),
	.OUT(n980));
   XOR2 U1708 (.A(n1548),
	.B(n1549),
	.OUT(n964));
   XOR2 U1709 (.A(n1551),
	.B(n2308),
	.OUT(n2307));
   XOR2 U1710 (.A(n1554),
	.B(n334),
	.OUT(n971));
   XOR2 U1711 (.A(n1556),
	.B(n1557),
	.OUT(n2309));
   XOR2 U1712 (.A(\mult_21/ab[4][5] ),
	.B(n329),
	.OUT(n983));
   XOR2 U1713 (.A(n1562),
	.B(n1563),
	.OUT(n2310));
   XOR2 U1714 (.A(n1565),
	.B(n341),
	.OUT(n986));
   XOR2 U1715 (.A(n1568),
	.B(n2311),
	.OUT(n989));
   XOR2 U1716 (.A(n1571),
	.B(n378),
	.OUT(n2312));
   XOR2 U1717 (.A(\mult_21/ab[7][3] ),
	.B(n380),
	.OUT(n991));
   XOR2 U1718 (.A(n343),
	.B(\mult_21/ab[2][2] ),
	.OUT(n994));
   XOR2 U1719 (.A(n1534),
	.B(n2314),
	.OUT(n2313));
   XOR2 U1720 (.A(\mult_21/ab[4][2] ),
	.B(n345),
	.OUT(n997));
   XOR2 U1721 (.A(n1546),
	.B(n2316),
	.OUT(n2315));
   XOR2 U1722 (.A(\mult_21/ab[6][2] ),
	.B(n347),
	.OUT(n1000));
   XOR2 U1723 (.A(\mult_21/ab[7][2] ),
	.B(n349),
	.OUT(n2317));
   XOR2 U1724 (.A(n351),
	.B(\mult_21/ab[2][1] ),
	.OUT(n1003));
   XOR2 U1725 (.A(n1578),
	.B(n2319),
	.OUT(n2318));
   XOR2 U1726 (.A(\mult_21/ab[4][1] ),
	.B(n353),
	.OUT(n1006));
   XOR2 U1727 (.A(n1583),
	.B(n1580),
	.OUT(n2320));
   XOR2 U1728 (.A(\mult_21/ab[6][1] ),
	.B(n355),
	.OUT(n1009));
   XOR2 U1729 (.A(\mult_21/ab[7][1] ),
	.B(n357),
	.OUT(n2321));
   XOR2 U1730 (.A(\mult_21/ab[6][5] ),
	.B(n373),
	.OUT(n1012));
   XOR2 U1731 (.A(\mult_21/ab[7][5] ),
	.B(n376),
	.OUT(n1014));
   XOR2 U1732 (.A(\mult_21/ab[7][4] ),
	.B(n2323),
	.OUT(n2322));
   XOR2 U1733 (.A(\mult_21/ab[7][0] ),
	.B(n365),
	.OUT(n1016));
   XOR2 U1734 (.A(n1600),
	.B(n363),
	.OUT(n2178));
   XOR2 U1735 (.A(n1597),
	.B(n1594),
	.OUT(n1017));
   XOR2 U1736 (.A(n1593),
	.B(n361),
	.OUT(n2179));
   XOR2 U1737 (.A(n1591),
	.B(n2324),
	.OUT(n1019));
   XOR2 U1738 (.A(n359),
	.B(\mult_21/ab[2][0] ),
	.OUT(n2180));
   XOR2 U1739 (.A(n1615),
	.B(\mult_20_3/ab[2][3] ),
	.OUT(n1034));
   XOR2 U1740 (.A(n1620),
	.B(\mult_20_3/ab[2][4] ),
	.OUT(n1031));
   XOR2 U1741 (.A(n1613),
	.B(n2326),
	.OUT(n2325));
   XOR2 U1742 (.A(n1630),
	.B(\mult_20_3/ab[2][5] ),
	.OUT(n1025));
   XOR2 U1743 (.A(n1618),
	.B(n2328),
	.OUT(n2327));
   XOR2 U1744 (.A(n1621),
	.B(n396),
	.OUT(n1037));
   XOR2 U1745 (.A(n1625),
	.B(n1626),
	.OUT(n1021));
   XOR2 U1746 (.A(n1628),
	.B(n2330),
	.OUT(n2329));
   XOR2 U1747 (.A(n1631),
	.B(n391),
	.OUT(n1028));
   XOR2 U1748 (.A(n1633),
	.B(n1634),
	.OUT(n2331));
   XOR2 U1749 (.A(\mult_20_3/ab[4][5] ),
	.B(n386),
	.OUT(n1040));
   XOR2 U1750 (.A(n1639),
	.B(n1640),
	.OUT(n2332));
   XOR2 U1751 (.A(n1642),
	.B(n398),
	.OUT(n1043));
   XOR2 U1752 (.A(n1645),
	.B(n2333),
	.OUT(n1046));
   XOR2 U1753 (.A(n1648),
	.B(n435),
	.OUT(n2334));
   XOR2 U1754 (.A(\mult_20_3/ab[7][3] ),
	.B(n437),
	.OUT(n1048));
   XOR2 U1755 (.A(n400),
	.B(\mult_20_3/ab[2][2] ),
	.OUT(n1051));
   XOR2 U1756 (.A(n1611),
	.B(n2336),
	.OUT(n2335));
   XOR2 U1757 (.A(\mult_20_3/ab[4][2] ),
	.B(n402),
	.OUT(n1054));
   XOR2 U1758 (.A(n1623),
	.B(n2338),
	.OUT(n2337));
   XOR2 U1759 (.A(\mult_20_3/ab[6][2] ),
	.B(n404),
	.OUT(n1057));
   XOR2 U1760 (.A(\mult_20_3/ab[7][2] ),
	.B(n406),
	.OUT(n2339));
   XOR2 U1761 (.A(n408),
	.B(\mult_20_3/ab[2][1] ),
	.OUT(n1060));
   XOR2 U1762 (.A(n1655),
	.B(n2341),
	.OUT(n2340));
   XOR2 U1763 (.A(\mult_20_3/ab[4][1] ),
	.B(n410),
	.OUT(n1063));
   XOR2 U1764 (.A(n1660),
	.B(n1657),
	.OUT(n2342));
   XOR2 U1765 (.A(\mult_20_3/ab[6][1] ),
	.B(n412),
	.OUT(n1066));
   XOR2 U1766 (.A(\mult_20_3/ab[7][1] ),
	.B(n414),
	.OUT(n2343));
   XOR2 U1767 (.A(\mult_20_3/ab[6][5] ),
	.B(n430),
	.OUT(n1069));
   XOR2 U1768 (.A(\mult_20_3/ab[7][5] ),
	.B(n433),
	.OUT(n1071));
   XOR2 U1769 (.A(\mult_20_3/ab[7][4] ),
	.B(n2345),
	.OUT(n2344));
   XOR2 U1770 (.A(\mult_20_3/ab[7][0] ),
	.B(n422),
	.OUT(n1073));
   XOR2 U1771 (.A(n1677),
	.B(n420),
	.OUT(n2181));
   XOR2 U1772 (.A(n1674),
	.B(n1671),
	.OUT(n1074));
   XOR2 U1773 (.A(n1670),
	.B(n418),
	.OUT(n2182));
   XOR2 U1774 (.A(n1668),
	.B(n2346),
	.OUT(n1076));
   XOR2 U1775 (.A(n416),
	.B(\mult_20_3/ab[2][0] ),
	.OUT(n2183));
   XOR2 U1776 (.A(n1692),
	.B(\mult_20_2/ab[2][3] ),
	.OUT(n1091));
   XOR2 U1777 (.A(n1697),
	.B(\mult_20_2/ab[2][4] ),
	.OUT(n1088));
   XOR2 U1778 (.A(n1690),
	.B(n2348),
	.OUT(n2347));
   XOR2 U1779 (.A(n1707),
	.B(\mult_20_2/ab[2][5] ),
	.OUT(n1082));
   XOR2 U1780 (.A(n1695),
	.B(n2350),
	.OUT(n2349));
   XOR2 U1781 (.A(n1698),
	.B(n453),
	.OUT(n1094));
   XOR2 U1782 (.A(n1702),
	.B(n1703),
	.OUT(n1078));
   XOR2 U1783 (.A(n1705),
	.B(n2352),
	.OUT(n2351));
   XOR2 U1784 (.A(n1708),
	.B(n448),
	.OUT(n1085));
   XOR2 U1785 (.A(n1710),
	.B(n1711),
	.OUT(n2353));
   XOR2 U1786 (.A(\mult_20_2/ab[4][5] ),
	.B(n443),
	.OUT(n1097));
   XOR2 U1787 (.A(n1716),
	.B(n1717),
	.OUT(n2354));
   XOR2 U1788 (.A(n1719),
	.B(n455),
	.OUT(n1100));
   XOR2 U1789 (.A(n1722),
	.B(n2355),
	.OUT(n1103));
   XOR2 U1790 (.A(n1725),
	.B(n492),
	.OUT(n2356));
   XOR2 U1791 (.A(\mult_20_2/ab[7][3] ),
	.B(n494),
	.OUT(n1105));
   XOR2 U1792 (.A(n457),
	.B(\mult_20_2/ab[2][2] ),
	.OUT(n1108));
   XOR2 U1793 (.A(n1688),
	.B(n2358),
	.OUT(n2357));
   XOR2 U1794 (.A(\mult_20_2/ab[4][2] ),
	.B(n459),
	.OUT(n1111));
   XOR2 U1795 (.A(n1700),
	.B(n2360),
	.OUT(n2359));
   XOR2 U1796 (.A(\mult_20_2/ab[6][2] ),
	.B(n461),
	.OUT(n1114));
   XOR2 U1797 (.A(\mult_20_2/ab[7][2] ),
	.B(n463),
	.OUT(n2361));
   XOR2 U1798 (.A(n465),
	.B(\mult_20_2/ab[2][1] ),
	.OUT(n1117));
   XOR2 U1799 (.A(n1732),
	.B(n2363),
	.OUT(n2362));
   XOR2 U1800 (.A(\mult_20_2/ab[4][1] ),
	.B(n467),
	.OUT(n1120));
   XOR2 U1801 (.A(n1737),
	.B(n1734),
	.OUT(n2364));
   XOR2 U1802 (.A(\mult_20_2/ab[6][1] ),
	.B(n469),
	.OUT(n1123));
   XOR2 U1803 (.A(\mult_20_2/ab[7][1] ),
	.B(n471),
	.OUT(n2365));
   XOR2 U1804 (.A(\mult_20_2/ab[6][5] ),
	.B(n487),
	.OUT(n1126));
   XOR2 U1805 (.A(\mult_20_2/ab[7][5] ),
	.B(n490),
	.OUT(n1128));
   XOR2 U1806 (.A(\mult_20_2/ab[7][4] ),
	.B(n2367),
	.OUT(n2366));
   XOR2 U1807 (.A(\mult_20_2/ab[7][0] ),
	.B(n479),
	.OUT(n1130));
   XOR2 U1808 (.A(n1754),
	.B(n477),
	.OUT(n2184));
   XOR2 U1809 (.A(n1751),
	.B(n1748),
	.OUT(n1131));
   XOR2 U1810 (.A(n1747),
	.B(n475),
	.OUT(n2185));
   XOR2 U1811 (.A(n1745),
	.B(n2368),
	.OUT(n1133));
   XOR2 U1812 (.A(n473),
	.B(\mult_20_2/ab[2][0] ),
	.OUT(n2186));
   XOR2 U1813 (.A(n1769),
	.B(\mult_20/ab[2][3] ),
	.OUT(n1148));
   XOR2 U1814 (.A(n1774),
	.B(\mult_20/ab[2][4] ),
	.OUT(n1145));
   XOR2 U1815 (.A(n1767),
	.B(n2370),
	.OUT(n2369));
   XOR2 U1816 (.A(n1784),
	.B(\mult_20/ab[2][5] ),
	.OUT(n1139));
   XOR2 U1817 (.A(n1772),
	.B(n2372),
	.OUT(n2371));
   XOR2 U1818 (.A(n1775),
	.B(n510),
	.OUT(n1151));
   XOR2 U1819 (.A(n1779),
	.B(n1780),
	.OUT(n1135));
   XOR2 U1820 (.A(n1782),
	.B(n2374),
	.OUT(n2373));
   XOR2 U1821 (.A(n1785),
	.B(n505),
	.OUT(n1142));
   XOR2 U1822 (.A(n1787),
	.B(n1788),
	.OUT(n2375));
   XOR2 U1823 (.A(\mult_20/ab[4][5] ),
	.B(n500),
	.OUT(n1154));
   XOR2 U1824 (.A(n1793),
	.B(n1794),
	.OUT(n2376));
   XOR2 U1825 (.A(n1796),
	.B(n512),
	.OUT(n1157));
   XOR2 U1826 (.A(n1799),
	.B(n2377),
	.OUT(n1160));
   XOR2 U1827 (.A(n1802),
	.B(n549),
	.OUT(n2378));
   XOR2 U1828 (.A(\mult_20/ab[7][3] ),
	.B(n551),
	.OUT(n1162));
   XOR2 U1829 (.A(n514),
	.B(\mult_20/ab[2][2] ),
	.OUT(n1165));
   XOR2 U1830 (.A(n1765),
	.B(n2380),
	.OUT(n2379));
   XOR2 U1831 (.A(\mult_20/ab[4][2] ),
	.B(n516),
	.OUT(n1168));
   XOR2 U1832 (.A(n1777),
	.B(n2382),
	.OUT(n2381));
   XOR2 U1833 (.A(\mult_20/ab[6][2] ),
	.B(n518),
	.OUT(n1171));
   XOR2 U1834 (.A(\mult_20/ab[7][2] ),
	.B(n520),
	.OUT(n2383));
   XOR2 U1835 (.A(n522),
	.B(\mult_20/ab[2][1] ),
	.OUT(n1174));
   XOR2 U1836 (.A(n1809),
	.B(n2385),
	.OUT(n2384));
   XOR2 U1837 (.A(\mult_20/ab[4][1] ),
	.B(n524),
	.OUT(n1177));
   XOR2 U1838 (.A(n1814),
	.B(n1811),
	.OUT(n2386));
   XOR2 U1839 (.A(\mult_20/ab[6][1] ),
	.B(n526),
	.OUT(n1180));
   XOR2 U1840 (.A(\mult_20/ab[7][1] ),
	.B(n528),
	.OUT(n2387));
   XOR2 U1841 (.A(\mult_20/ab[6][5] ),
	.B(n544),
	.OUT(n1183));
   XOR2 U1842 (.A(\mult_20/ab[7][5] ),
	.B(n547),
	.OUT(n1185));
   XOR2 U1843 (.A(\mult_20/ab[7][4] ),
	.B(n2389),
	.OUT(n2388));
   XOR2 U1844 (.A(\mult_20/ab[7][0] ),
	.B(n536),
	.OUT(n1187));
   XOR2 U1845 (.A(n1831),
	.B(n534),
	.OUT(n2187));
   XOR2 U1846 (.A(n1828),
	.B(n1825),
	.OUT(n1188));
   XOR2 U1847 (.A(n1824),
	.B(n532),
	.OUT(n2188));
   XOR2 U1848 (.A(n1822),
	.B(n2390),
	.OUT(n1190));
   XOR2 U1849 (.A(n530),
	.B(\mult_20/ab[2][0] ),
	.OUT(n2189));
   XOR2 U1850 (.A(n1846),
	.B(\mult_19_3/ab[2][3] ),
	.OUT(n1205));
   XOR2 U1851 (.A(n1851),
	.B(\mult_19_3/ab[2][4] ),
	.OUT(n1202));
   XOR2 U1852 (.A(n1844),
	.B(n2392),
	.OUT(n2391));
   XOR2 U1853 (.A(n1861),
	.B(\mult_19_3/ab[2][5] ),
	.OUT(n1196));
   XOR2 U1854 (.A(n1849),
	.B(n2394),
	.OUT(n2393));
   XOR2 U1855 (.A(n1852),
	.B(n567),
	.OUT(n1208));
   XOR2 U1856 (.A(n1856),
	.B(n1857),
	.OUT(n1192));
   XOR2 U1857 (.A(n1859),
	.B(n2396),
	.OUT(n2395));
   XOR2 U1858 (.A(n1862),
	.B(n562),
	.OUT(n1199));
   XOR2 U1859 (.A(n1864),
	.B(n1865),
	.OUT(n2397));
   XOR2 U1860 (.A(\mult_19_3/ab[4][5] ),
	.B(n557),
	.OUT(n1211));
   XOR2 U1861 (.A(n1870),
	.B(n1871),
	.OUT(n2398));
   XOR2 U1862 (.A(n1873),
	.B(n569),
	.OUT(n1214));
   XOR2 U1863 (.A(n1876),
	.B(n2399),
	.OUT(n1217));
   XOR2 U1864 (.A(n1879),
	.B(n606),
	.OUT(n2400));
   XOR2 U1865 (.A(\mult_19_3/ab[7][3] ),
	.B(n608),
	.OUT(n1219));
   XOR2 U1866 (.A(n571),
	.B(\mult_19_3/ab[2][2] ),
	.OUT(n1222));
   XOR2 U1867 (.A(n1842),
	.B(n2402),
	.OUT(n2401));
   XOR2 U1868 (.A(\mult_19_3/ab[4][2] ),
	.B(n573),
	.OUT(n1225));
   XOR2 U1869 (.A(n1854),
	.B(n2404),
	.OUT(n2403));
   XOR2 U1870 (.A(\mult_19_3/ab[6][2] ),
	.B(n575),
	.OUT(n1228));
   XOR2 U1871 (.A(\mult_19_3/ab[7][2] ),
	.B(n577),
	.OUT(n2405));
   XOR2 U1872 (.A(n579),
	.B(\mult_19_3/ab[2][1] ),
	.OUT(n1231));
   XOR2 U1873 (.A(n1886),
	.B(n2407),
	.OUT(n2406));
   XOR2 U1874 (.A(\mult_19_3/ab[4][1] ),
	.B(n581),
	.OUT(n1234));
   XOR2 U1875 (.A(n1891),
	.B(n1888),
	.OUT(n2408));
   XOR2 U1876 (.A(\mult_19_3/ab[6][1] ),
	.B(n583),
	.OUT(n1237));
   XOR2 U1877 (.A(\mult_19_3/ab[7][1] ),
	.B(n585),
	.OUT(n2409));
   XOR2 U1878 (.A(\mult_19_3/ab[6][5] ),
	.B(n601),
	.OUT(n1240));
   XOR2 U1879 (.A(\mult_19_3/ab[7][5] ),
	.B(n604),
	.OUT(n1242));
   XOR2 U1880 (.A(\mult_19_3/ab[7][4] ),
	.B(n2411),
	.OUT(n2410));
   XOR2 U1881 (.A(\mult_19_3/ab[7][0] ),
	.B(n593),
	.OUT(n1244));
   XOR2 U1882 (.A(n1908),
	.B(n591),
	.OUT(n2190));
   XOR2 U1883 (.A(n1905),
	.B(n1902),
	.OUT(n1245));
   XOR2 U1884 (.A(n1901),
	.B(n589),
	.OUT(n2191));
   XOR2 U1885 (.A(n1899),
	.B(n2412),
	.OUT(n1247));
   XOR2 U1886 (.A(n587),
	.B(\mult_19_3/ab[2][0] ),
	.OUT(n2192));
   XOR2 U1887 (.A(n1923),
	.B(\mult_19_2/ab[2][3] ),
	.OUT(n1262));
   XOR2 U1888 (.A(n1928),
	.B(\mult_19_2/ab[2][4] ),
	.OUT(n1259));
   XOR2 U1889 (.A(n1921),
	.B(n2414),
	.OUT(n2413));
   XOR2 U1890 (.A(n1938),
	.B(\mult_19_2/ab[2][5] ),
	.OUT(n1253));
   XOR2 U1891 (.A(n1926),
	.B(n2416),
	.OUT(n2415));
   XOR2 U1892 (.A(n1929),
	.B(n624),
	.OUT(n1265));
   XOR2 U1893 (.A(n1933),
	.B(n1934),
	.OUT(n1249));
   XOR2 U1894 (.A(n1936),
	.B(n2418),
	.OUT(n2417));
   XOR2 U1895 (.A(n1939),
	.B(n619),
	.OUT(n1256));
   XOR2 U1896 (.A(n1941),
	.B(n1942),
	.OUT(n2419));
   XOR2 U1897 (.A(\mult_19_2/ab[4][5] ),
	.B(n614),
	.OUT(n1268));
   XOR2 U1898 (.A(n1947),
	.B(n1948),
	.OUT(n2420));
   XOR2 U1899 (.A(n1950),
	.B(n626),
	.OUT(n1271));
   XOR2 U1900 (.A(n1953),
	.B(n2421),
	.OUT(n1274));
   XOR2 U1901 (.A(n1956),
	.B(n663),
	.OUT(n2422));
   XOR2 U1902 (.A(\mult_19_2/ab[7][3] ),
	.B(n665),
	.OUT(n1276));
   XOR2 U1903 (.A(n628),
	.B(\mult_19_2/ab[2][2] ),
	.OUT(n1279));
   XOR2 U1904 (.A(n1919),
	.B(n2424),
	.OUT(n2423));
   XOR2 U1905 (.A(\mult_19_2/ab[4][2] ),
	.B(n630),
	.OUT(n1282));
   XOR2 U1906 (.A(n1931),
	.B(n2426),
	.OUT(n2425));
   XOR2 U1907 (.A(\mult_19_2/ab[6][2] ),
	.B(n632),
	.OUT(n1285));
   XOR2 U1908 (.A(\mult_19_2/ab[7][2] ),
	.B(n634),
	.OUT(n2427));
   XOR2 U1909 (.A(n636),
	.B(\mult_19_2/ab[2][1] ),
	.OUT(n1288));
   XOR2 U1910 (.A(n1963),
	.B(n2429),
	.OUT(n2428));
   XOR2 U1911 (.A(\mult_19_2/ab[4][1] ),
	.B(n638),
	.OUT(n1291));
   XOR2 U1912 (.A(n1968),
	.B(n1965),
	.OUT(n2430));
   XOR2 U1913 (.A(\mult_19_2/ab[6][1] ),
	.B(n640),
	.OUT(n1294));
   XOR2 U1914 (.A(\mult_19_2/ab[7][1] ),
	.B(n642),
	.OUT(n2431));
   XOR2 U1915 (.A(\mult_19_2/ab[6][5] ),
	.B(n658),
	.OUT(n1297));
   XOR2 U1916 (.A(\mult_19_2/ab[7][5] ),
	.B(n661),
	.OUT(n1299));
   XOR2 U1917 (.A(\mult_19_2/ab[7][4] ),
	.B(n2433),
	.OUT(n2432));
   XOR2 U1918 (.A(\mult_19_2/ab[7][0] ),
	.B(n650),
	.OUT(n1301));
   XOR2 U1919 (.A(n1985),
	.B(n648),
	.OUT(n2193));
   XOR2 U1920 (.A(n1982),
	.B(n1979),
	.OUT(n1302));
   XOR2 U1921 (.A(n1978),
	.B(n646),
	.OUT(n2194));
   XOR2 U1922 (.A(n1976),
	.B(n2434),
	.OUT(n1304));
   XOR2 U1923 (.A(n644),
	.B(\mult_19_2/ab[2][0] ),
	.OUT(n2195));
   XOR2 U1924 (.A(n2000),
	.B(\mult_19/ab[2][3] ),
	.OUT(n1319));
   XOR2 U1925 (.A(n2005),
	.B(\mult_19/ab[2][4] ),
	.OUT(n1316));
   XOR2 U1926 (.A(n1998),
	.B(n2436),
	.OUT(n2435));
   XOR2 U1927 (.A(n2015),
	.B(\mult_19/ab[2][5] ),
	.OUT(n1310));
   XOR2 U1928 (.A(n2003),
	.B(n2438),
	.OUT(n2437));
   XOR2 U1929 (.A(n2006),
	.B(n681),
	.OUT(n1322));
   XOR2 U1930 (.A(n2010),
	.B(n2011),
	.OUT(n1306));
   XOR2 U1931 (.A(n2013),
	.B(n2440),
	.OUT(n2439));
   XOR2 U1932 (.A(n2016),
	.B(n676),
	.OUT(n1313));
   XOR2 U1933 (.A(n2018),
	.B(n2019),
	.OUT(n2441));
   XOR2 U1934 (.A(\mult_19/ab[4][5] ),
	.B(n671),
	.OUT(n1325));
   XOR2 U1935 (.A(n2024),
	.B(n2025),
	.OUT(n2442));
   XOR2 U1936 (.A(n2027),
	.B(n683),
	.OUT(n1328));
   XOR2 U1937 (.A(n2030),
	.B(n2443),
	.OUT(n1331));
   XOR2 U1938 (.A(n2033),
	.B(n720),
	.OUT(n2444));
   XOR2 U1939 (.A(\mult_19/ab[7][3] ),
	.B(n722),
	.OUT(n1333));
   XOR2 U1940 (.A(n685),
	.B(\mult_19/ab[2][2] ),
	.OUT(n1336));
   XOR2 U1941 (.A(n1996),
	.B(n2446),
	.OUT(n2445));
   XOR2 U1942 (.A(\mult_19/ab[4][2] ),
	.B(n687),
	.OUT(n1339));
   XOR2 U1943 (.A(n2008),
	.B(n2448),
	.OUT(n2447));
   XOR2 U1944 (.A(\mult_19/ab[6][2] ),
	.B(n689),
	.OUT(n1342));
   XOR2 U1945 (.A(\mult_19/ab[7][2] ),
	.B(n691),
	.OUT(n2449));
   XOR2 U1946 (.A(n693),
	.B(\mult_19/ab[2][1] ),
	.OUT(n1345));
   XOR2 U1947 (.A(n2040),
	.B(n2451),
	.OUT(n2450));
   XOR2 U1948 (.A(\mult_19/ab[4][1] ),
	.B(n695),
	.OUT(n1348));
   XOR2 U1949 (.A(n2045),
	.B(n2042),
	.OUT(n2452));
   XOR2 U1950 (.A(\mult_19/ab[6][1] ),
	.B(n697),
	.OUT(n1351));
   XOR2 U1951 (.A(\mult_19/ab[7][1] ),
	.B(n699),
	.OUT(n2453));
   XOR2 U1952 (.A(\mult_19/ab[6][5] ),
	.B(n715),
	.OUT(n1354));
   XOR2 U1953 (.A(\mult_19/ab[7][5] ),
	.B(n718),
	.OUT(n1356));
   XOR2 U1954 (.A(\mult_19/ab[7][4] ),
	.B(n2455),
	.OUT(n2454));
   XOR2 U1955 (.A(\mult_19/ab[7][0] ),
	.B(n707),
	.OUT(n1358));
   XOR2 U1956 (.A(n2062),
	.B(n705),
	.OUT(n2196));
   XOR2 U1957 (.A(n2059),
	.B(n2056),
	.OUT(n1359));
   XOR2 U1958 (.A(n2055),
	.B(n703),
	.OUT(n2197));
   XOR2 U1959 (.A(n2053),
	.B(n2456),
	.OUT(n1361));
   XOR2 U1960 (.A(n701),
	.B(\mult_19/ab[2][0] ),
	.OUT(n2198));
   XOR2 U1961 (.A(n2070),
	.B(n2457),
	.OUT(n1366));
   XOR2 U1962 (.A(N3),
	.B(N19),
	.OUT(n2458));
   XOR2 U1963 (.A(N16),
	.B(N32),
	.OUT(n2459));
   XOR2 U1964 (.A(N64),
	.B(n2459),
	.OUT(n2199));
   XOR2 U1965 (.A(n2460),
	.B(n2461),
	.OUT(n2200));
   XOR2 U1966 (.A(N63),
	.B(n2462),
	.OUT(n2202));
   XOR2 U1967 (.A(N62),
	.B(n762),
	.OUT(n2203));
   XOR2 U1968 (.A(N61),
	.B(n759),
	.OUT(n2204));
   XOR2 U1969 (.A(N60),
	.B(n757),
	.OUT(n2205));
   XOR2 U1970 (.A(N59),
	.B(n754),
	.OUT(n2206));
   XOR2 U1971 (.A(N58),
	.B(n752),
	.OUT(n2207));
   XOR2 U1972 (.A(N57),
	.B(n749),
	.OUT(n2208));
   XOR2 U1973 (.A(N56),
	.B(n2089),
	.OUT(n2209));
   XOR2 U1974 (.A(N55),
	.B(n2086),
	.OUT(n2211));
   XOR2 U1975 (.A(N54),
	.B(n745),
	.OUT(n2212));
   XOR2 U1976 (.A(N53),
	.B(n742),
	.OUT(n2213));
   XOR2 U1977 (.A(N52),
	.B(n2075),
	.OUT(n2215));
   XOR2 U1978 (.A(n739),
	.B(n2076),
	.OUT(n2217));
   XOR2 U1979 (.A(n736),
	.B(n737),
	.OUT(n2218));
   XOR2 U1980 (.A(n2104),
	.B(n2463),
	.OUT(n1371));
   XOR2 U1981 (.A(N163),
	.B(N179),
	.OUT(n2464));
   XOR2 U1982 (.A(N176),
	.B(N192),
	.OUT(n2465));
   XOR2 U1983 (.A(N224),
	.B(n2465),
	.OUT(n2219));
   XOR2 U1984 (.A(n2466),
	.B(n2467),
	.OUT(n2220));
   XOR2 U1985 (.A(N223),
	.B(n2468),
	.OUT(n2222));
   XOR2 U1986 (.A(N222),
	.B(n804),
	.OUT(n2223));
   XOR2 U1987 (.A(N221),
	.B(n801),
	.OUT(n2224));
   XOR2 U1988 (.A(N220),
	.B(n799),
	.OUT(n2225));
   XOR2 U1989 (.A(N219),
	.B(n796),
	.OUT(n2226));
   XOR2 U1990 (.A(N218),
	.B(n794),
	.OUT(n2227));
   XOR2 U1991 (.A(N217),
	.B(n791),
	.OUT(n2228));
   XOR2 U1992 (.A(N216),
	.B(n2123),
	.OUT(n2229));
   XOR2 U1993 (.A(N215),
	.B(n2120),
	.OUT(n2231));
   XOR2 U1994 (.A(N214),
	.B(n787),
	.OUT(n2232));
   XOR2 U1995 (.A(N213),
	.B(n784),
	.OUT(n2233));
   XOR2 U1996 (.A(N212),
	.B(n2109),
	.OUT(n2235));
   XOR2 U1997 (.A(n781),
	.B(n2110),
	.OUT(n2237));
   XOR2 U1998 (.A(n778),
	.B(n779),
	.OUT(n2238));
   XOR2 U1999 (.A(n2138),
	.B(n2469),
	.OUT(n1376));
   XOR2 U2000 (.A(N83),
	.B(N99),
	.OUT(n2470));
   XOR2 U2001 (.A(N96),
	.B(N112),
	.OUT(n2471));
   XOR2 U2002 (.A(N144),
	.B(n2471),
	.OUT(n2239));
   XOR2 U2003 (.A(n2472),
	.B(n2473),
	.OUT(n2240));
   XOR2 U2004 (.A(N143),
	.B(n2474),
	.OUT(n2242));
   XOR2 U2005 (.A(N142),
	.B(n846),
	.OUT(n2243));
   XOR2 U2006 (.A(N141),
	.B(n843),
	.OUT(n2244));
   XOR2 U2007 (.A(N140),
	.B(n841),
	.OUT(n2245));
   XOR2 U2008 (.A(N139),
	.B(n838),
	.OUT(n2246));
   XOR2 U2009 (.A(N138),
	.B(n836),
	.OUT(n2247));
   XOR2 U2010 (.A(N137),
	.B(n833),
	.OUT(n2248));
   XOR2 U2011 (.A(N136),
	.B(n2157),
	.OUT(n2249));
   XOR2 U2012 (.A(N135),
	.B(n2154),
	.OUT(n2251));
   XOR2 U2013 (.A(N134),
	.B(n829),
	.OUT(n2252));
   XOR2 U2014 (.A(N133),
	.B(n826),
	.OUT(n2253));
   XOR2 U2015 (.A(N132),
	.B(n2143),
	.OUT(n2255));
   XOR2 U2016 (.A(n823),
	.B(n2144),
	.OUT(n2257));
   XOR2 U2017 (.A(n820),
	.B(n821),
	.OUT(n2258));
   INVERTER U2018 (.IN(n669),
	.OUT(n2015));
   INVERTER U2019 (.IN(n674),
	.OUT(n2005));
   INVERTER U2020 (.IN(n679),
	.OUT(n2000));
   INVERTER U2021 (.IN(n612),
	.OUT(n1938));
   INVERTER U2022 (.IN(n617),
	.OUT(n1928));
   INVERTER U2023 (.IN(n622),
	.OUT(n1923));
   INVERTER U2024 (.IN(n2070),
	.OUT(n2475));
   INVERTER U2025 (.IN(n555),
	.OUT(n1861));
   INVERTER U2026 (.IN(n560),
	.OUT(n1851));
   INVERTER U2027 (.IN(n565),
	.OUT(n1846));
   INVERTER U2028 (.IN(n498),
	.OUT(n1784));
   INVERTER U2029 (.IN(n503),
	.OUT(n1774));
   INVERTER U2030 (.IN(n508),
	.OUT(n1769));
   INVERTER U2031 (.IN(n441),
	.OUT(n1707));
   INVERTER U2032 (.IN(n446),
	.OUT(n1697));
   INVERTER U2033 (.IN(n451),
	.OUT(n1692));
   INVERTER U2034 (.IN(n2138),
	.OUT(n2476));
   INVERTER U2035 (.IN(n384),
	.OUT(n1630));
   INVERTER U2036 (.IN(n389),
	.OUT(n1620));
   INVERTER U2037 (.IN(n394),
	.OUT(n1615));
   INVERTER U2038 (.IN(n327),
	.OUT(n1553));
   INVERTER U2039 (.IN(n332),
	.OUT(n1543));
   INVERTER U2040 (.IN(n337),
	.OUT(n1538));
   INVERTER U2041 (.IN(n270),
	.OUT(n1476));
   INVERTER U2042 (.IN(n275),
	.OUT(n1466));
   INVERTER U2043 (.IN(n280),
	.OUT(n1461));
   INVERTER U2044 (.IN(n2104),
	.OUT(n2477));
   INVERTER U2045 (.IN(n213),
	.OUT(n1399));
   INVERTER U2046 (.IN(n218),
	.OUT(n1389));
   INVERTER U2047 (.IN(n223),
	.OUT(n1384));
   OAI22 U2048 (.OUT(n2478),
	.D(n1394),
	.C(n1396),
	.B(n210),
	.A(n1395));
   OAI21 U2049 (.OUT(n2479),
	.C(n2478),
	.B(\mult_21_3/ab[3][6] ),
	.A(\mult_21_3/ab[2][7] ));
   OAI21 U2050 (.OUT(n2480),
	.C(n2479),
	.B(n2482),
	.A(n2481));
   INVERTER U2051 (.IN(n1398),
	.OUT(n2264));
   OAI21 U2052 (.OUT(n1407),
	.C(n849),
	.B(n2264),
	.A(\mult_21_3/ab[3][5] ));
   INVERTER U2053 (.IN(n1415),
	.OUT(n2267));
   INVERTER U2054 (.IN(n1388),
	.OUT(n2262));
   OAI21 U2055 (.OUT(n1401),
	.C(n853),
	.B(n2262),
	.A(\mult_21_3/ab[3][4] ));
   INVERTER U2056 (.IN(n220),
	.OUT(n1410));
   INVERTER U2057 (.IN(n1409),
	.OUT(n1418));
   OAI21 U2058 (.OUT(n1419),
	.C(n867),
	.B(n1409),
	.A(\mult_21_3/ab[5][4] ));
   INVERTER U2059 (.IN(n264),
	.OUT(n1452));
   INVERTER U2060 (.IN(n1383),
	.OUT(n2260));
   OAI21 U2061 (.OUT(n1391),
	.C(n859),
	.B(n2260),
	.A(\mult_21_3/ab[3][3] ));
   INVERTER U2062 (.IN(n225),
	.OUT(n1404));
   INVERTER U2063 (.IN(n1403),
	.OUT(n1412));
   OAI21 U2064 (.OUT(n1413),
	.C(n855),
	.B(n1403),
	.A(\mult_21_3/ab[5][3] ));
   INVERTER U2065 (.IN(n227),
	.OUT(n1420));
   INVERTER U2066 (.IN(n1378),
	.OUT(n2270));
   OAI21 U2067 (.OUT(n1381),
	.C(n862),
	.B(n2270),
	.A(\mult_21_3/ab[3][2] ));
   INVERTER U2068 (.IN(n1385),
	.OUT(n2272));
   OAI21 U2069 (.OUT(n1393),
	.C(n864),
	.B(n2272),
	.A(\mult_21_3/ab[5][2] ));
   AOI22 U2070 (.A(n235),
	.B(\mult_21_3/ab[7][2] ),
	.C(n2483),
	.D(n870),
	.OUT(n204));
   INVERTER U2071 (.IN(n1422),
	.OUT(n2275));
   OAI21 U2072 (.OUT(n1425),
	.C(n879),
	.B(n2275),
	.A(\mult_21_3/ab[3][1] ));
   INVERTER U2073 (.IN(n1426),
	.OUT(n1430));
   OAI21 U2074 (.OUT(n1431),
	.C(n881),
	.B(n1426),
	.A(\mult_21_3/ab[5][1] ));
   AOI22 U2075 (.A(n243),
	.B(\mult_21_3/ab[7][1] ),
	.C(n2484),
	.D(n2485),
	.OUT(n206));
   INVERTER U2076 (.IN(n1435),
	.OUT(n2280));
   OAI21 U2077 (.OUT(n1438),
	.C(n888),
	.B(n2280),
	.A(\mult_21_3/ab[3][0] ));
   INVERTER U2078 (.IN(n247),
	.OUT(n1441));
   INVERTER U2079 (.IN(n1440),
	.OUT(n1444));
   OAI21 U2080 (.OUT(n1445),
	.C(n2486),
	.B(n1440),
	.A(\mult_21_3/ab[5][0] ));
   INVERTER U2081 (.IN(n249),
	.OUT(n1447));
   AOI22 U2082 (.A(n251),
	.B(\mult_21_3/ab[7][0] ),
	.C(n2487),
	.D(n901),
	.OUT(n208));
   AOI22 U2083 (.A(\mult_21_3/ab[4][6] ),
	.B(\mult_21_3/ab[3][7] ),
	.C(n2480),
	.D(n2489),
	.OUT(n2488));
   OAI22 U2084 (.OUT(n2490),
	.D(n253),
	.C(n2492),
	.B(n2488),
	.A(n2491));
   AOI22 U2085 (.A(\mult_21_3/ab[5][7] ),
	.B(\mult_21_3/ab[6][6] ),
	.C(n2490),
	.D(n254),
	.OUT(n2493));
   AOI22 U2086 (.A(\mult_21_3/ab[6][7] ),
	.B(\mult_21_3/ab[7][6] ),
	.C(n2494),
	.D(n2495),
	.OUT(n194));
   OAI21 U2087 (.OUT(n1449),
	.C(n874),
	.B(n2267),
	.A(\mult_21_3/ab[5][5] ));
   OAI22 U2088 (.OUT(n197),
	.D(n899),
	.C(n261),
	.B(n2496),
	.A(n262));
   INVERTER U2089 (.IN(n1451),
	.OUT(n2279));
   OAI21 U2090 (.OUT(n2497),
	.C(n896),
	.B(n1451),
	.A(\mult_21_3/ab[7][4] ));
   OAI21 U2091 (.OUT(n200),
	.C(n2497),
	.B(n1453),
	.A(n2279));
   AOI22 U2092 (.A(n266),
	.B(\mult_21_3/ab[7][3] ),
	.C(n2498),
	.D(n2499),
	.OUT(n202));
   OAI22 U2093 (.OUT(n2500),
	.D(n1471),
	.C(n1473),
	.B(n267),
	.A(n1472));
   OAI21 U2094 (.OUT(n2501),
	.C(n2500),
	.B(\mult_21_2/ab[3][6] ),
	.A(\mult_21_2/ab[2][7] ));
   OAI21 U2095 (.OUT(n2502),
	.C(n2501),
	.B(n2504),
	.A(n2503));
   INVERTER U2096 (.IN(n1475),
	.OUT(n2286));
   OAI21 U2097 (.OUT(n1484),
	.C(n906),
	.B(n2286),
	.A(\mult_21_2/ab[3][5] ));
   INVERTER U2098 (.IN(n1492),
	.OUT(n2289));
   INVERTER U2099 (.IN(n1465),
	.OUT(n2284));
   OAI21 U2100 (.OUT(n1478),
	.C(n910),
	.B(n2284),
	.A(\mult_21_2/ab[3][4] ));
   INVERTER U2101 (.IN(n277),
	.OUT(n1487));
   INVERTER U2102 (.IN(n1486),
	.OUT(n1495));
   OAI21 U2103 (.OUT(n1496),
	.C(n924),
	.B(n1486),
	.A(\mult_21_2/ab[5][4] ));
   INVERTER U2104 (.IN(n321),
	.OUT(n1529));
   INVERTER U2105 (.IN(n1460),
	.OUT(n2282));
   OAI21 U2106 (.OUT(n1468),
	.C(n916),
	.B(n2282),
	.A(\mult_21_2/ab[3][3] ));
   INVERTER U2107 (.IN(n282),
	.OUT(n1481));
   INVERTER U2108 (.IN(n1480),
	.OUT(n1489));
   OAI21 U2109 (.OUT(n1490),
	.C(n912),
	.B(n1480),
	.A(\mult_21_2/ab[5][3] ));
   INVERTER U2110 (.IN(n284),
	.OUT(n1497));
   INVERTER U2111 (.IN(n1455),
	.OUT(n2292));
   OAI21 U2112 (.OUT(n1458),
	.C(n919),
	.B(n2292),
	.A(\mult_21_2/ab[3][2] ));
   INVERTER U2113 (.IN(n1462),
	.OUT(n2294));
   OAI21 U2114 (.OUT(n1470),
	.C(n921),
	.B(n2294),
	.A(\mult_21_2/ab[5][2] ));
   AOI22 U2115 (.A(n292),
	.B(\mult_21_2/ab[7][2] ),
	.C(n2505),
	.D(n927),
	.OUT(n188));
   INVERTER U2116 (.IN(n1499),
	.OUT(n2297));
   OAI21 U2117 (.OUT(n1502),
	.C(n936),
	.B(n2297),
	.A(\mult_21_2/ab[3][1] ));
   INVERTER U2118 (.IN(n1503),
	.OUT(n1507));
   OAI21 U2119 (.OUT(n1508),
	.C(n938),
	.B(n1503),
	.A(\mult_21_2/ab[5][1] ));
   AOI22 U2120 (.A(n300),
	.B(\mult_21_2/ab[7][1] ),
	.C(n2506),
	.D(n2507),
	.OUT(n190));
   INVERTER U2121 (.IN(n1512),
	.OUT(n2302));
   OAI21 U2122 (.OUT(n1515),
	.C(n945),
	.B(n2302),
	.A(\mult_21_2/ab[3][0] ));
   INVERTER U2123 (.IN(n304),
	.OUT(n1518));
   INVERTER U2124 (.IN(n1517),
	.OUT(n1521));
   OAI21 U2125 (.OUT(n1522),
	.C(n2508),
	.B(n1517),
	.A(\mult_21_2/ab[5][0] ));
   INVERTER U2126 (.IN(n306),
	.OUT(n1524));
   AOI22 U2127 (.A(n308),
	.B(\mult_21_2/ab[7][0] ),
	.C(n2509),
	.D(n958),
	.OUT(n192));
   AOI22 U2128 (.A(\mult_21_2/ab[4][6] ),
	.B(\mult_21_2/ab[3][7] ),
	.C(n2502),
	.D(n2511),
	.OUT(n2510));
   OAI22 U2129 (.OUT(n2512),
	.D(n310),
	.C(n2514),
	.B(n2510),
	.A(n2513));
   AOI22 U2130 (.A(\mult_21_2/ab[5][7] ),
	.B(\mult_21_2/ab[6][6] ),
	.C(n2512),
	.D(n311),
	.OUT(n2515));
   AOI22 U2131 (.A(\mult_21_2/ab[6][7] ),
	.B(\mult_21_2/ab[7][6] ),
	.C(n2516),
	.D(n2517),
	.OUT(n178));
   OAI21 U2132 (.OUT(n1526),
	.C(n931),
	.B(n2289),
	.A(\mult_21_2/ab[5][5] ));
   OAI22 U2133 (.OUT(n181),
	.D(n956),
	.C(n318),
	.B(n2518),
	.A(n319));
   INVERTER U2134 (.IN(n1528),
	.OUT(n2301));
   OAI21 U2135 (.OUT(n2519),
	.C(n953),
	.B(n1528),
	.A(\mult_21_2/ab[7][4] ));
   OAI21 U2136 (.OUT(n184),
	.C(n2519),
	.B(n1530),
	.A(n2301));
   AOI22 U2137 (.A(n323),
	.B(\mult_21_2/ab[7][3] ),
	.C(n2520),
	.D(n2521),
	.OUT(n186));
   OAI22 U2138 (.OUT(n2522),
	.D(n1548),
	.C(n1550),
	.B(n324),
	.A(n1549));
   OAI21 U2139 (.OUT(n2523),
	.C(n2522),
	.B(\mult_21/ab[3][6] ),
	.A(\mult_21/ab[2][7] ));
   OAI21 U2140 (.OUT(n2524),
	.C(n2523),
	.B(n2526),
	.A(n2525));
   INVERTER U2141 (.IN(n1552),
	.OUT(n2308));
   OAI21 U2142 (.OUT(n1561),
	.C(n963),
	.B(n2308),
	.A(\mult_21/ab[3][5] ));
   INVERTER U2143 (.IN(n1569),
	.OUT(n2311));
   INVERTER U2144 (.IN(n1542),
	.OUT(n2306));
   OAI21 U2145 (.OUT(n1555),
	.C(n967),
	.B(n2306),
	.A(\mult_21/ab[3][4] ));
   INVERTER U2146 (.IN(n334),
	.OUT(n1564));
   INVERTER U2147 (.IN(n1563),
	.OUT(n1572));
   OAI21 U2148 (.OUT(n1573),
	.C(n981),
	.B(n1563),
	.A(\mult_21/ab[5][4] ));
   INVERTER U2149 (.IN(n378),
	.OUT(n1606));
   INVERTER U2150 (.IN(n1537),
	.OUT(n2304));
   OAI21 U2151 (.OUT(n1545),
	.C(n973),
	.B(n2304),
	.A(\mult_21/ab[3][3] ));
   INVERTER U2152 (.IN(n339),
	.OUT(n1558));
   INVERTER U2153 (.IN(n1557),
	.OUT(n1566));
   OAI21 U2154 (.OUT(n1567),
	.C(n969),
	.B(n1557),
	.A(\mult_21/ab[5][3] ));
   INVERTER U2155 (.IN(n341),
	.OUT(n1574));
   INVERTER U2156 (.IN(n1532),
	.OUT(n2314));
   OAI21 U2157 (.OUT(n1535),
	.C(n976),
	.B(n2314),
	.A(\mult_21/ab[3][2] ));
   INVERTER U2158 (.IN(n1539),
	.OUT(n2316));
   OAI21 U2159 (.OUT(n1547),
	.C(n978),
	.B(n2316),
	.A(\mult_21/ab[5][2] ));
   AOI22 U2160 (.A(n349),
	.B(\mult_21/ab[7][2] ),
	.C(n2527),
	.D(n984),
	.OUT(n172));
   INVERTER U2161 (.IN(n1576),
	.OUT(n2319));
   OAI21 U2162 (.OUT(n1579),
	.C(n993),
	.B(n2319),
	.A(\mult_21/ab[3][1] ));
   INVERTER U2163 (.IN(n1580),
	.OUT(n1584));
   OAI21 U2164 (.OUT(n1585),
	.C(n995),
	.B(n1580),
	.A(\mult_21/ab[5][1] ));
   AOI22 U2165 (.A(n357),
	.B(\mult_21/ab[7][1] ),
	.C(n2528),
	.D(n2529),
	.OUT(n174));
   INVERTER U2166 (.IN(n1589),
	.OUT(n2324));
   OAI21 U2167 (.OUT(n1592),
	.C(n1002),
	.B(n2324),
	.A(\mult_21/ab[3][0] ));
   INVERTER U2168 (.IN(n361),
	.OUT(n1595));
   INVERTER U2169 (.IN(n1594),
	.OUT(n1598));
   OAI21 U2170 (.OUT(n1599),
	.C(n2530),
	.B(n1594),
	.A(\mult_21/ab[5][0] ));
   INVERTER U2171 (.IN(n363),
	.OUT(n1601));
   AOI22 U2172 (.A(n365),
	.B(\mult_21/ab[7][0] ),
	.C(n2531),
	.D(n1015),
	.OUT(n176));
   AOI22 U2173 (.A(\mult_21/ab[4][6] ),
	.B(\mult_21/ab[3][7] ),
	.C(n2524),
	.D(n2533),
	.OUT(n2532));
   OAI22 U2174 (.OUT(n2534),
	.D(n367),
	.C(n2536),
	.B(n2532),
	.A(n2535));
   AOI22 U2175 (.A(\mult_21/ab[5][7] ),
	.B(\mult_21/ab[6][6] ),
	.C(n2534),
	.D(n368),
	.OUT(n2537));
   AOI22 U2176 (.A(\mult_21/ab[6][7] ),
	.B(\mult_21/ab[7][6] ),
	.C(n2538),
	.D(n2539),
	.OUT(n162));
   OAI21 U2177 (.OUT(n1603),
	.C(n988),
	.B(n2311),
	.A(\mult_21/ab[5][5] ));
   OAI22 U2178 (.OUT(n165),
	.D(n1013),
	.C(n375),
	.B(n2540),
	.A(n376));
   INVERTER U2179 (.IN(n1605),
	.OUT(n2323));
   OAI21 U2180 (.OUT(n2541),
	.C(n1010),
	.B(n1605),
	.A(\mult_21/ab[7][4] ));
   OAI21 U2181 (.OUT(n168),
	.C(n2541),
	.B(n1607),
	.A(n2323));
   AOI22 U2182 (.A(n380),
	.B(\mult_21/ab[7][3] ),
	.C(n2542),
	.D(n2543),
	.OUT(n170));
   OAI22 U2183 (.OUT(n2544),
	.D(n1625),
	.C(n1627),
	.B(n381),
	.A(n1626));
   OAI21 U2184 (.OUT(n2545),
	.C(n2544),
	.B(\mult_20_3/ab[3][6] ),
	.A(\mult_20_3/ab[2][7] ));
   OAI21 U2185 (.OUT(n2546),
	.C(n2545),
	.B(n2548),
	.A(n2547));
   INVERTER U2186 (.IN(n1629),
	.OUT(n2330));
   OAI21 U2187 (.OUT(n1638),
	.C(n1020),
	.B(n2330),
	.A(\mult_20_3/ab[3][5] ));
   INVERTER U2188 (.IN(n1646),
	.OUT(n2333));
   INVERTER U2189 (.IN(n1619),
	.OUT(n2328));
   OAI21 U2190 (.OUT(n1632),
	.C(n1024),
	.B(n2328),
	.A(\mult_20_3/ab[3][4] ));
   INVERTER U2191 (.IN(n391),
	.OUT(n1641));
   INVERTER U2192 (.IN(n1640),
	.OUT(n1649));
   OAI21 U2193 (.OUT(n1650),
	.C(n1038),
	.B(n1640),
	.A(\mult_20_3/ab[5][4] ));
   INVERTER U2194 (.IN(n435),
	.OUT(n1683));
   INVERTER U2195 (.IN(n1614),
	.OUT(n2326));
   OAI21 U2196 (.OUT(n1622),
	.C(n1030),
	.B(n2326),
	.A(\mult_20_3/ab[3][3] ));
   INVERTER U2197 (.IN(n396),
	.OUT(n1635));
   INVERTER U2198 (.IN(n1634),
	.OUT(n1643));
   OAI21 U2199 (.OUT(n1644),
	.C(n1026),
	.B(n1634),
	.A(\mult_20_3/ab[5][3] ));
   INVERTER U2200 (.IN(n398),
	.OUT(n1651));
   INVERTER U2201 (.IN(n1609),
	.OUT(n2336));
   OAI21 U2202 (.OUT(n1612),
	.C(n1033),
	.B(n2336),
	.A(\mult_20_3/ab[3][2] ));
   INVERTER U2203 (.IN(n1616),
	.OUT(n2338));
   OAI21 U2204 (.OUT(n1624),
	.C(n1035),
	.B(n2338),
	.A(\mult_20_3/ab[5][2] ));
   AOI22 U2205 (.A(n406),
	.B(\mult_20_3/ab[7][2] ),
	.C(n2549),
	.D(n1041),
	.OUT(n156));
   INVERTER U2206 (.IN(n1653),
	.OUT(n2341));
   OAI21 U2207 (.OUT(n1656),
	.C(n1050),
	.B(n2341),
	.A(\mult_20_3/ab[3][1] ));
   INVERTER U2208 (.IN(n1657),
	.OUT(n1661));
   OAI21 U2209 (.OUT(n1662),
	.C(n1052),
	.B(n1657),
	.A(\mult_20_3/ab[5][1] ));
   AOI22 U2210 (.A(n414),
	.B(\mult_20_3/ab[7][1] ),
	.C(n2550),
	.D(n2551),
	.OUT(n158));
   INVERTER U2211 (.IN(n1666),
	.OUT(n2346));
   OAI21 U2212 (.OUT(n1669),
	.C(n1059),
	.B(n2346),
	.A(\mult_20_3/ab[3][0] ));
   INVERTER U2213 (.IN(n418),
	.OUT(n1672));
   INVERTER U2214 (.IN(n1671),
	.OUT(n1675));
   OAI21 U2215 (.OUT(n1676),
	.C(n2552),
	.B(n1671),
	.A(\mult_20_3/ab[5][0] ));
   INVERTER U2216 (.IN(n420),
	.OUT(n1678));
   AOI22 U2217 (.A(n422),
	.B(\mult_20_3/ab[7][0] ),
	.C(n2553),
	.D(n1072),
	.OUT(n160));
   AOI22 U2218 (.A(\mult_20_3/ab[4][6] ),
	.B(\mult_20_3/ab[3][7] ),
	.C(n2546),
	.D(n2555),
	.OUT(n2554));
   OAI22 U2219 (.OUT(n2556),
	.D(n424),
	.C(n2558),
	.B(n2554),
	.A(n2557));
   AOI22 U2220 (.A(\mult_20_3/ab[5][7] ),
	.B(\mult_20_3/ab[6][6] ),
	.C(n2556),
	.D(n425),
	.OUT(n2559));
   AOI22 U2221 (.A(\mult_20_3/ab[6][7] ),
	.B(\mult_20_3/ab[7][6] ),
	.C(n2560),
	.D(n2561),
	.OUT(n146));
   OAI21 U2222 (.OUT(n1680),
	.C(n1045),
	.B(n2333),
	.A(\mult_20_3/ab[5][5] ));
   OAI22 U2223 (.OUT(n149),
	.D(n1070),
	.C(n432),
	.B(n2562),
	.A(n433));
   INVERTER U2224 (.IN(n1682),
	.OUT(n2345));
   OAI21 U2225 (.OUT(n2563),
	.C(n1067),
	.B(n1682),
	.A(\mult_20_3/ab[7][4] ));
   OAI21 U2226 (.OUT(n152),
	.C(n2563),
	.B(n1684),
	.A(n2345));
   AOI22 U2227 (.A(n437),
	.B(\mult_20_3/ab[7][3] ),
	.C(n2564),
	.D(n2565),
	.OUT(n154));
   OAI22 U2228 (.OUT(n2566),
	.D(n1702),
	.C(n1704),
	.B(n438),
	.A(n1703));
   OAI21 U2229 (.OUT(n2567),
	.C(n2566),
	.B(\mult_20_2/ab[3][6] ),
	.A(\mult_20_2/ab[2][7] ));
   OAI21 U2230 (.OUT(n2568),
	.C(n2567),
	.B(n2570),
	.A(n2569));
   INVERTER U2231 (.IN(n1706),
	.OUT(n2352));
   OAI21 U2232 (.OUT(n1715),
	.C(n1077),
	.B(n2352),
	.A(\mult_20_2/ab[3][5] ));
   INVERTER U2233 (.IN(n1723),
	.OUT(n2355));
   INVERTER U2234 (.IN(n1696),
	.OUT(n2350));
   OAI21 U2235 (.OUT(n1709),
	.C(n1081),
	.B(n2350),
	.A(\mult_20_2/ab[3][4] ));
   INVERTER U2236 (.IN(n448),
	.OUT(n1718));
   INVERTER U2237 (.IN(n1717),
	.OUT(n1726));
   OAI21 U2238 (.OUT(n1727),
	.C(n1095),
	.B(n1717),
	.A(\mult_20_2/ab[5][4] ));
   INVERTER U2239 (.IN(n492),
	.OUT(n1760));
   INVERTER U2240 (.IN(n1691),
	.OUT(n2348));
   OAI21 U2241 (.OUT(n1699),
	.C(n1087),
	.B(n2348),
	.A(\mult_20_2/ab[3][3] ));
   INVERTER U2242 (.IN(n453),
	.OUT(n1712));
   INVERTER U2243 (.IN(n1711),
	.OUT(n1720));
   OAI21 U2244 (.OUT(n1721),
	.C(n1083),
	.B(n1711),
	.A(\mult_20_2/ab[5][3] ));
   INVERTER U2245 (.IN(n455),
	.OUT(n1728));
   INVERTER U2246 (.IN(n1686),
	.OUT(n2358));
   OAI21 U2247 (.OUT(n1689),
	.C(n1090),
	.B(n2358),
	.A(\mult_20_2/ab[3][2] ));
   INVERTER U2248 (.IN(n1693),
	.OUT(n2360));
   OAI21 U2249 (.OUT(n1701),
	.C(n1092),
	.B(n2360),
	.A(\mult_20_2/ab[5][2] ));
   AOI22 U2250 (.A(n463),
	.B(\mult_20_2/ab[7][2] ),
	.C(n2571),
	.D(n1098),
	.OUT(n140));
   INVERTER U2251 (.IN(n1730),
	.OUT(n2363));
   OAI21 U2252 (.OUT(n1733),
	.C(n1107),
	.B(n2363),
	.A(\mult_20_2/ab[3][1] ));
   INVERTER U2253 (.IN(n1734),
	.OUT(n1738));
   OAI21 U2254 (.OUT(n1739),
	.C(n1109),
	.B(n1734),
	.A(\mult_20_2/ab[5][1] ));
   AOI22 U2255 (.A(n471),
	.B(\mult_20_2/ab[7][1] ),
	.C(n2572),
	.D(n2573),
	.OUT(n142));
   INVERTER U2256 (.IN(n1743),
	.OUT(n2368));
   OAI21 U2257 (.OUT(n1746),
	.C(n1116),
	.B(n2368),
	.A(\mult_20_2/ab[3][0] ));
   INVERTER U2258 (.IN(n475),
	.OUT(n1749));
   INVERTER U2259 (.IN(n1748),
	.OUT(n1752));
   OAI21 U2260 (.OUT(n1753),
	.C(n2574),
	.B(n1748),
	.A(\mult_20_2/ab[5][0] ));
   INVERTER U2261 (.IN(n477),
	.OUT(n1755));
   AOI22 U2262 (.A(n479),
	.B(\mult_20_2/ab[7][0] ),
	.C(n2575),
	.D(n1129),
	.OUT(n144));
   AOI22 U2263 (.A(\mult_20_2/ab[4][6] ),
	.B(\mult_20_2/ab[3][7] ),
	.C(n2568),
	.D(n2577),
	.OUT(n2576));
   OAI22 U2264 (.OUT(n2578),
	.D(n481),
	.C(n2580),
	.B(n2576),
	.A(n2579));
   AOI22 U2265 (.A(\mult_20_2/ab[5][7] ),
	.B(\mult_20_2/ab[6][6] ),
	.C(n2578),
	.D(n482),
	.OUT(n2581));
   AOI22 U2266 (.A(\mult_20_2/ab[6][7] ),
	.B(\mult_20_2/ab[7][6] ),
	.C(n2582),
	.D(n2583),
	.OUT(n130));
   OAI21 U2267 (.OUT(n1757),
	.C(n1102),
	.B(n2355),
	.A(\mult_20_2/ab[5][5] ));
   OAI22 U2268 (.OUT(n133),
	.D(n1127),
	.C(n489),
	.B(n2584),
	.A(n490));
   INVERTER U2269 (.IN(n1759),
	.OUT(n2367));
   OAI21 U2270 (.OUT(n2585),
	.C(n1124),
	.B(n1759),
	.A(\mult_20_2/ab[7][4] ));
   OAI21 U2271 (.OUT(n136),
	.C(n2585),
	.B(n1761),
	.A(n2367));
   AOI22 U2272 (.A(n494),
	.B(\mult_20_2/ab[7][3] ),
	.C(n2586),
	.D(n2587),
	.OUT(n138));
   OAI22 U2273 (.OUT(n2588),
	.D(n1779),
	.C(n1781),
	.B(n495),
	.A(n1780));
   OAI21 U2274 (.OUT(n2589),
	.C(n2588),
	.B(\mult_20/ab[3][6] ),
	.A(\mult_20/ab[2][7] ));
   OAI21 U2275 (.OUT(n2590),
	.C(n2589),
	.B(n2592),
	.A(n2591));
   INVERTER U2276 (.IN(n1783),
	.OUT(n2374));
   OAI21 U2277 (.OUT(n1792),
	.C(n1134),
	.B(n2374),
	.A(\mult_20/ab[3][5] ));
   INVERTER U2278 (.IN(n1800),
	.OUT(n2377));
   INVERTER U2279 (.IN(n1773),
	.OUT(n2372));
   OAI21 U2280 (.OUT(n1786),
	.C(n1138),
	.B(n2372),
	.A(\mult_20/ab[3][4] ));
   INVERTER U2281 (.IN(n505),
	.OUT(n1795));
   INVERTER U2282 (.IN(n1794),
	.OUT(n1803));
   OAI21 U2283 (.OUT(n1804),
	.C(n1152),
	.B(n1794),
	.A(\mult_20/ab[5][4] ));
   INVERTER U2284 (.IN(n549),
	.OUT(n1837));
   INVERTER U2285 (.IN(n1768),
	.OUT(n2370));
   OAI21 U2286 (.OUT(n1776),
	.C(n1144),
	.B(n2370),
	.A(\mult_20/ab[3][3] ));
   INVERTER U2287 (.IN(n510),
	.OUT(n1789));
   INVERTER U2288 (.IN(n1788),
	.OUT(n1797));
   OAI21 U2289 (.OUT(n1798),
	.C(n1140),
	.B(n1788),
	.A(\mult_20/ab[5][3] ));
   INVERTER U2290 (.IN(n512),
	.OUT(n1805));
   INVERTER U2291 (.IN(n1763),
	.OUT(n2380));
   OAI21 U2292 (.OUT(n1766),
	.C(n1147),
	.B(n2380),
	.A(\mult_20/ab[3][2] ));
   INVERTER U2293 (.IN(n1770),
	.OUT(n2382));
   OAI21 U2294 (.OUT(n1778),
	.C(n1149),
	.B(n2382),
	.A(\mult_20/ab[5][2] ));
   AOI22 U2295 (.A(n520),
	.B(\mult_20/ab[7][2] ),
	.C(n2593),
	.D(n1155),
	.OUT(n124));
   INVERTER U2296 (.IN(n1807),
	.OUT(n2385));
   OAI21 U2297 (.OUT(n1810),
	.C(n1164),
	.B(n2385),
	.A(\mult_20/ab[3][1] ));
   INVERTER U2298 (.IN(n1811),
	.OUT(n1815));
   OAI21 U2299 (.OUT(n1816),
	.C(n1166),
	.B(n1811),
	.A(\mult_20/ab[5][1] ));
   AOI22 U2300 (.A(n528),
	.B(\mult_20/ab[7][1] ),
	.C(n2594),
	.D(n2595),
	.OUT(n126));
   INVERTER U2301 (.IN(n1820),
	.OUT(n2390));
   OAI21 U2302 (.OUT(n1823),
	.C(n1173),
	.B(n2390),
	.A(\mult_20/ab[3][0] ));
   INVERTER U2303 (.IN(n532),
	.OUT(n1826));
   INVERTER U2304 (.IN(n1825),
	.OUT(n1829));
   OAI21 U2305 (.OUT(n1830),
	.C(n2596),
	.B(n1825),
	.A(\mult_20/ab[5][0] ));
   INVERTER U2306 (.IN(n534),
	.OUT(n1832));
   AOI22 U2307 (.A(n536),
	.B(\mult_20/ab[7][0] ),
	.C(n2597),
	.D(n1186),
	.OUT(n128));
   AOI22 U2308 (.A(\mult_20/ab[4][6] ),
	.B(\mult_20/ab[3][7] ),
	.C(n2590),
	.D(n2599),
	.OUT(n2598));
   OAI22 U2309 (.OUT(n2600),
	.D(n538),
	.C(n2602),
	.B(n2598),
	.A(n2601));
   AOI22 U2310 (.A(\mult_20/ab[5][7] ),
	.B(\mult_20/ab[6][6] ),
	.C(n2600),
	.D(n539),
	.OUT(n2603));
   AOI22 U2311 (.A(\mult_20/ab[6][7] ),
	.B(\mult_20/ab[7][6] ),
	.C(n2604),
	.D(n2605),
	.OUT(n114));
   OAI21 U2312 (.OUT(n1834),
	.C(n1159),
	.B(n2377),
	.A(\mult_20/ab[5][5] ));
   OAI22 U2313 (.OUT(n117),
	.D(n1184),
	.C(n546),
	.B(n2606),
	.A(n547));
   INVERTER U2314 (.IN(n1836),
	.OUT(n2389));
   OAI21 U2315 (.OUT(n2607),
	.C(n1181),
	.B(n1836),
	.A(\mult_20/ab[7][4] ));
   OAI21 U2316 (.OUT(n120),
	.C(n2607),
	.B(n1838),
	.A(n2389));
   AOI22 U2317 (.A(n551),
	.B(\mult_20/ab[7][3] ),
	.C(n2608),
	.D(n2609),
	.OUT(n122));
   OAI22 U2318 (.OUT(n2610),
	.D(n1856),
	.C(n1858),
	.B(n552),
	.A(n1857));
   OAI21 U2319 (.OUT(n2611),
	.C(n2610),
	.B(\mult_19_3/ab[3][6] ),
	.A(\mult_19_3/ab[2][7] ));
   OAI21 U2320 (.OUT(n2612),
	.C(n2611),
	.B(n2614),
	.A(n2613));
   INVERTER U2321 (.IN(n1860),
	.OUT(n2396));
   OAI21 U2322 (.OUT(n1869),
	.C(n1191),
	.B(n2396),
	.A(\mult_19_3/ab[3][5] ));
   INVERTER U2323 (.IN(n1877),
	.OUT(n2399));
   INVERTER U2324 (.IN(n1850),
	.OUT(n2394));
   OAI21 U2325 (.OUT(n1863),
	.C(n1195),
	.B(n2394),
	.A(\mult_19_3/ab[3][4] ));
   INVERTER U2326 (.IN(n562),
	.OUT(n1872));
   INVERTER U2327 (.IN(n1871),
	.OUT(n1880));
   OAI21 U2328 (.OUT(n1881),
	.C(n1209),
	.B(n1871),
	.A(\mult_19_3/ab[5][4] ));
   INVERTER U2329 (.IN(n606),
	.OUT(n1914));
   INVERTER U2330 (.IN(n1845),
	.OUT(n2392));
   OAI21 U2331 (.OUT(n1853),
	.C(n1201),
	.B(n2392),
	.A(\mult_19_3/ab[3][3] ));
   INVERTER U2332 (.IN(n567),
	.OUT(n1866));
   INVERTER U2333 (.IN(n1865),
	.OUT(n1874));
   OAI21 U2334 (.OUT(n1875),
	.C(n1197),
	.B(n1865),
	.A(\mult_19_3/ab[5][3] ));
   INVERTER U2335 (.IN(n569),
	.OUT(n1882));
   INVERTER U2336 (.IN(n1840),
	.OUT(n2402));
   OAI21 U2337 (.OUT(n1843),
	.C(n1204),
	.B(n2402),
	.A(\mult_19_3/ab[3][2] ));
   INVERTER U2338 (.IN(n1847),
	.OUT(n2404));
   OAI21 U2339 (.OUT(n1855),
	.C(n1206),
	.B(n2404),
	.A(\mult_19_3/ab[5][2] ));
   AOI22 U2340 (.A(n577),
	.B(\mult_19_3/ab[7][2] ),
	.C(n2615),
	.D(n1212),
	.OUT(n108));
   INVERTER U2341 (.IN(n1884),
	.OUT(n2407));
   OAI21 U2342 (.OUT(n1887),
	.C(n1221),
	.B(n2407),
	.A(\mult_19_3/ab[3][1] ));
   INVERTER U2343 (.IN(n1888),
	.OUT(n1892));
   OAI21 U2344 (.OUT(n1893),
	.C(n1223),
	.B(n1888),
	.A(\mult_19_3/ab[5][1] ));
   AOI22 U2345 (.A(n585),
	.B(\mult_19_3/ab[7][1] ),
	.C(n2616),
	.D(n2617),
	.OUT(n110));
   INVERTER U2346 (.IN(n1897),
	.OUT(n2412));
   OAI21 U2347 (.OUT(n1900),
	.C(n1230),
	.B(n2412),
	.A(\mult_19_3/ab[3][0] ));
   INVERTER U2348 (.IN(n589),
	.OUT(n1903));
   INVERTER U2349 (.IN(n1902),
	.OUT(n1906));
   OAI21 U2350 (.OUT(n1907),
	.C(n2618),
	.B(n1902),
	.A(\mult_19_3/ab[5][0] ));
   INVERTER U2351 (.IN(n591),
	.OUT(n1909));
   AOI22 U2352 (.A(n593),
	.B(\mult_19_3/ab[7][0] ),
	.C(n2619),
	.D(n1243),
	.OUT(n112));
   AOI22 U2353 (.A(\mult_19_3/ab[4][6] ),
	.B(\mult_19_3/ab[3][7] ),
	.C(n2612),
	.D(n2621),
	.OUT(n2620));
   OAI22 U2354 (.OUT(n2622),
	.D(n595),
	.C(n2624),
	.B(n2620),
	.A(n2623));
   AOI22 U2355 (.A(\mult_19_3/ab[5][7] ),
	.B(\mult_19_3/ab[6][6] ),
	.C(n2622),
	.D(n596),
	.OUT(n2625));
   AOI22 U2356 (.A(\mult_19_3/ab[6][7] ),
	.B(\mult_19_3/ab[7][6] ),
	.C(n2626),
	.D(n2627),
	.OUT(n98));
   OAI21 U2357 (.OUT(n1911),
	.C(n1216),
	.B(n2399),
	.A(\mult_19_3/ab[5][5] ));
   OAI22 U2358 (.OUT(n101),
	.D(n1241),
	.C(n603),
	.B(n2628),
	.A(n604));
   INVERTER U2359 (.IN(n1913),
	.OUT(n2411));
   OAI21 U2360 (.OUT(n2629),
	.C(n1238),
	.B(n1913),
	.A(\mult_19_3/ab[7][4] ));
   OAI21 U2361 (.OUT(n104),
	.C(n2629),
	.B(n1915),
	.A(n2411));
   AOI22 U2362 (.A(n608),
	.B(\mult_19_3/ab[7][3] ),
	.C(n2630),
	.D(n2631),
	.OUT(n106));
   OAI22 U2363 (.OUT(n2632),
	.D(n1933),
	.C(n1935),
	.B(n609),
	.A(n1934));
   OAI21 U2364 (.OUT(n2633),
	.C(n2632),
	.B(\mult_19_2/ab[3][6] ),
	.A(\mult_19_2/ab[2][7] ));
   OAI21 U2365 (.OUT(n2634),
	.C(n2633),
	.B(n2636),
	.A(n2635));
   INVERTER U2366 (.IN(n1937),
	.OUT(n2418));
   OAI21 U2367 (.OUT(n1946),
	.C(n1248),
	.B(n2418),
	.A(\mult_19_2/ab[3][5] ));
   INVERTER U2368 (.IN(n1954),
	.OUT(n2421));
   INVERTER U2369 (.IN(n1927),
	.OUT(n2416));
   OAI21 U2370 (.OUT(n1940),
	.C(n1252),
	.B(n2416),
	.A(\mult_19_2/ab[3][4] ));
   INVERTER U2371 (.IN(n619),
	.OUT(n1949));
   INVERTER U2372 (.IN(n1948),
	.OUT(n1957));
   OAI21 U2373 (.OUT(n1958),
	.C(n1266),
	.B(n1948),
	.A(\mult_19_2/ab[5][4] ));
   INVERTER U2374 (.IN(n663),
	.OUT(n1991));
   INVERTER U2375 (.IN(n1922),
	.OUT(n2414));
   OAI21 U2376 (.OUT(n1930),
	.C(n1258),
	.B(n2414),
	.A(\mult_19_2/ab[3][3] ));
   INVERTER U2377 (.IN(n624),
	.OUT(n1943));
   INVERTER U2378 (.IN(n1942),
	.OUT(n1951));
   OAI21 U2379 (.OUT(n1952),
	.C(n1254),
	.B(n1942),
	.A(\mult_19_2/ab[5][3] ));
   INVERTER U2380 (.IN(n626),
	.OUT(n1959));
   INVERTER U2381 (.IN(n1917),
	.OUT(n2424));
   OAI21 U2382 (.OUT(n1920),
	.C(n1261),
	.B(n2424),
	.A(\mult_19_2/ab[3][2] ));
   INVERTER U2383 (.IN(n1924),
	.OUT(n2426));
   OAI21 U2384 (.OUT(n1932),
	.C(n1263),
	.B(n2426),
	.A(\mult_19_2/ab[5][2] ));
   AOI22 U2385 (.A(n634),
	.B(\mult_19_2/ab[7][2] ),
	.C(n2637),
	.D(n1269),
	.OUT(n92));
   INVERTER U2386 (.IN(n1961),
	.OUT(n2429));
   OAI21 U2387 (.OUT(n1964),
	.C(n1278),
	.B(n2429),
	.A(\mult_19_2/ab[3][1] ));
   INVERTER U2388 (.IN(n1965),
	.OUT(n1969));
   OAI21 U2389 (.OUT(n1970),
	.C(n1280),
	.B(n1965),
	.A(\mult_19_2/ab[5][1] ));
   AOI22 U2390 (.A(n642),
	.B(\mult_19_2/ab[7][1] ),
	.C(n2638),
	.D(n2639),
	.OUT(n94));
   INVERTER U2391 (.IN(n1974),
	.OUT(n2434));
   OAI21 U2392 (.OUT(n1977),
	.C(n1287),
	.B(n2434),
	.A(\mult_19_2/ab[3][0] ));
   INVERTER U2393 (.IN(n646),
	.OUT(n1980));
   INVERTER U2394 (.IN(n1979),
	.OUT(n1983));
   OAI21 U2395 (.OUT(n1984),
	.C(n2640),
	.B(n1979),
	.A(\mult_19_2/ab[5][0] ));
   INVERTER U2396 (.IN(n648),
	.OUT(n1986));
   AOI22 U2397 (.A(n650),
	.B(\mult_19_2/ab[7][0] ),
	.C(n2641),
	.D(n1300),
	.OUT(n96));
   AOI22 U2398 (.A(\mult_19_2/ab[4][6] ),
	.B(\mult_19_2/ab[3][7] ),
	.C(n2634),
	.D(n2643),
	.OUT(n2642));
   OAI22 U2399 (.OUT(n2644),
	.D(n652),
	.C(n2646),
	.B(n2642),
	.A(n2645));
   AOI22 U2400 (.A(\mult_19_2/ab[5][7] ),
	.B(\mult_19_2/ab[6][6] ),
	.C(n2644),
	.D(n653),
	.OUT(n2647));
   AOI22 U2401 (.A(\mult_19_2/ab[6][7] ),
	.B(\mult_19_2/ab[7][6] ),
	.C(n2648),
	.D(n2649),
	.OUT(n82));
   OAI21 U2402 (.OUT(n1988),
	.C(n1273),
	.B(n2421),
	.A(\mult_19_2/ab[5][5] ));
   OAI22 U2403 (.OUT(n85),
	.D(n1298),
	.C(n660),
	.B(n2650),
	.A(n661));
   INVERTER U2404 (.IN(n1990),
	.OUT(n2433));
   OAI21 U2405 (.OUT(n2651),
	.C(n1295),
	.B(n1990),
	.A(\mult_19_2/ab[7][4] ));
   OAI21 U2406 (.OUT(n88),
	.C(n2651),
	.B(n1992),
	.A(n2433));
   AOI22 U2407 (.A(n665),
	.B(\mult_19_2/ab[7][3] ),
	.C(n2652),
	.D(n2653),
	.OUT(n90));
   OAI22 U2408 (.OUT(n2654),
	.D(n2010),
	.C(n2012),
	.B(n666),
	.A(n2011));
   OAI21 U2409 (.OUT(n2655),
	.C(n2654),
	.B(\mult_19/ab[3][6] ),
	.A(\mult_19/ab[2][7] ));
   OAI21 U2410 (.OUT(n2656),
	.C(n2655),
	.B(n2658),
	.A(n2657));
   INVERTER U2411 (.IN(n2014),
	.OUT(n2440));
   OAI21 U2412 (.OUT(n2023),
	.C(n1305),
	.B(n2440),
	.A(\mult_19/ab[3][5] ));
   INVERTER U2413 (.IN(n2031),
	.OUT(n2443));
   INVERTER U2414 (.IN(n2004),
	.OUT(n2438));
   OAI21 U2415 (.OUT(n2017),
	.C(n1309),
	.B(n2438),
	.A(\mult_19/ab[3][4] ));
   INVERTER U2416 (.IN(n676),
	.OUT(n2026));
   INVERTER U2417 (.IN(n2025),
	.OUT(n2034));
   OAI21 U2418 (.OUT(n2035),
	.C(n1323),
	.B(n2025),
	.A(\mult_19/ab[5][4] ));
   INVERTER U2419 (.IN(n720),
	.OUT(n2068));
   INVERTER U2420 (.IN(n1999),
	.OUT(n2436));
   OAI21 U2421 (.OUT(n2007),
	.C(n1315),
	.B(n2436),
	.A(\mult_19/ab[3][3] ));
   INVERTER U2422 (.IN(n681),
	.OUT(n2020));
   INVERTER U2423 (.IN(n2019),
	.OUT(n2028));
   OAI21 U2424 (.OUT(n2029),
	.C(n1311),
	.B(n2019),
	.A(\mult_19/ab[5][3] ));
   INVERTER U2425 (.IN(n683),
	.OUT(n2036));
   INVERTER U2426 (.IN(n1994),
	.OUT(n2446));
   OAI21 U2427 (.OUT(n1997),
	.C(n1318),
	.B(n2446),
	.A(\mult_19/ab[3][2] ));
   INVERTER U2428 (.IN(n2001),
	.OUT(n2448));
   OAI21 U2429 (.OUT(n2009),
	.C(n1320),
	.B(n2448),
	.A(\mult_19/ab[5][2] ));
   AOI22 U2430 (.A(n691),
	.B(\mult_19/ab[7][2] ),
	.C(n2659),
	.D(n1326),
	.OUT(n76));
   INVERTER U2431 (.IN(n2038),
	.OUT(n2451));
   OAI21 U2432 (.OUT(n2041),
	.C(n1335),
	.B(n2451),
	.A(\mult_19/ab[3][1] ));
   INVERTER U2433 (.IN(n2042),
	.OUT(n2046));
   OAI21 U2434 (.OUT(n2047),
	.C(n1337),
	.B(n2042),
	.A(\mult_19/ab[5][1] ));
   AOI22 U2435 (.A(n699),
	.B(\mult_19/ab[7][1] ),
	.C(n2660),
	.D(n2661),
	.OUT(n78));
   INVERTER U2436 (.IN(n2051),
	.OUT(n2456));
   OAI21 U2437 (.OUT(n2054),
	.C(n1344),
	.B(n2456),
	.A(\mult_19/ab[3][0] ));
   INVERTER U2438 (.IN(n703),
	.OUT(n2057));
   INVERTER U2439 (.IN(n2056),
	.OUT(n2060));
   OAI21 U2440 (.OUT(n2061),
	.C(n2662),
	.B(n2056),
	.A(\mult_19/ab[5][0] ));
   INVERTER U2441 (.IN(n705),
	.OUT(n2063));
   AOI22 U2442 (.A(n707),
	.B(\mult_19/ab[7][0] ),
	.C(n2663),
	.D(n1357),
	.OUT(n80));
   AOI22 U2443 (.A(\mult_19/ab[4][6] ),
	.B(\mult_19/ab[3][7] ),
	.C(n2656),
	.D(n2665),
	.OUT(n2664));
   OAI22 U2444 (.OUT(n2666),
	.D(n709),
	.C(n2668),
	.B(n2664),
	.A(n2667));
   AOI22 U2445 (.A(\mult_19/ab[5][7] ),
	.B(\mult_19/ab[6][6] ),
	.C(n2666),
	.D(n710),
	.OUT(n2669));
   AOI22 U2446 (.A(\mult_19/ab[6][7] ),
	.B(\mult_19/ab[7][6] ),
	.C(n2670),
	.D(n2671),
	.OUT(n66));
   OAI21 U2447 (.OUT(n2065),
	.C(n1330),
	.B(n2443),
	.A(\mult_19/ab[5][5] ));
   OAI22 U2448 (.OUT(n69),
	.D(n1355),
	.C(n717),
	.B(n2672),
	.A(n718));
   INVERTER U2449 (.IN(n2067),
	.OUT(n2455));
   OAI21 U2450 (.OUT(n2673),
	.C(n1352),
	.B(n2067),
	.A(\mult_19/ab[7][4] ));
   OAI21 U2451 (.OUT(n72),
	.C(n2673),
	.B(n2069),
	.A(n2455));
   AOI22 U2452 (.A(n722),
	.B(\mult_19/ab[7][3] ),
	.C(n2674),
	.D(n2675),
	.OUT(n74));
   OAI21 U2453 (.OUT(n2676),
	.C(n1363),
	.B(n1362),
	.A(n2475));
   OAI21 U2454 (.OUT(n2677),
	.C(n2676),
	.B(n2070),
	.A(n2457));
   OAI21 U2455 (.OUT(n2678),
	.C(n2677),
	.B(N3),
	.A(N19));
   AOI21 U2456 (.OUT(n2679),
	.C(n2680),
	.B(N3),
	.A(N19));
   OAI22 U2457 (.OUT(n2681),
	.D(n723),
	.C(n2683),
	.B(n2679),
	.A(n2682));
   AOI22 U2458 (.A(N21),
	.B(N5),
	.C(n2681),
	.D(n2685),
	.OUT(n2684));
   OAI22 U2459 (.OUT(n2686),
	.D(n725),
	.C(n2688),
	.B(n2684),
	.A(n2687));
   AOI22 U2460 (.A(N23),
	.B(N7),
	.C(n2686),
	.D(n2690),
	.OUT(n2689));
   OAI22 U2461 (.OUT(n2691),
	.D(n727),
	.C(n2693),
	.B(n2689),
	.A(n2692));
   AOI22 U2462 (.A(N25),
	.B(N9),
	.C(n2691),
	.D(n2695),
	.OUT(n2694));
   OAI22 U2463 (.OUT(n2696),
	.D(n729),
	.C(n2698),
	.B(n2694),
	.A(n2697));
   AOI22 U2464 (.A(N27),
	.B(N11),
	.C(n2696),
	.D(n2700),
	.OUT(n2699));
   OAI22 U2465 (.OUT(n2701),
	.D(n731),
	.C(n2703),
	.B(n2699),
	.A(n2702));
   AOI22 U2466 (.A(N29),
	.B(N13),
	.C(n2701),
	.D(n2705),
	.OUT(n2704));
   AOI22 U2467 (.A(N30),
	.B(N14),
	.C(n2707),
	.D(n2708),
	.OUT(n2706));
   OAI22 U2468 (.OUT(n2460),
	.D(n734),
	.C(n2072),
	.B(n2706),
	.A(n2071));
   AOI21 U2469 (.OUT(n2709),
	.C(n2214),
	.B(n2075),
	.A(n2078));
   INVERTER U2470 (.IN(n2082),
	.OUT(n2086));
   OAI21 U2471 (.OUT(n2087),
	.C(n2710),
	.B(n2082),
	.A(N55));
   INVERTER U2472 (.IN(n747),
	.OUT(n2089));
   INVERTER U2473 (.IN(n764),
	.OUT(n2462));
   OAI22 U2474 (.OUT(n2461),
	.D(n2201),
	.C(n2103),
	.B(n763),
	.A(n2462));
   OAI21 U2475 (.OUT(n2711),
	.C(n1368),
	.B(n1367),
	.A(n2477));
   OAI21 U2476 (.OUT(n2712),
	.C(n2711),
	.B(n2104),
	.A(n2463));
   OAI21 U2477 (.OUT(n2713),
	.C(n2712),
	.B(N163),
	.A(N179));
   AOI21 U2478 (.OUT(n2714),
	.C(n2715),
	.B(N163),
	.A(N179));
   OAI22 U2479 (.OUT(n2716),
	.D(n765),
	.C(n2718),
	.B(n2714),
	.A(n2717));
   AOI22 U2480 (.A(N181),
	.B(N165),
	.C(n2716),
	.D(n2720),
	.OUT(n2719));
   OAI22 U2481 (.OUT(n2721),
	.D(n767),
	.C(n2723),
	.B(n2719),
	.A(n2722));
   AOI22 U2482 (.A(N183),
	.B(N167),
	.C(n2721),
	.D(n2725),
	.OUT(n2724));
   OAI22 U2483 (.OUT(n2726),
	.D(n769),
	.C(n2728),
	.B(n2724),
	.A(n2727));
   AOI22 U2484 (.A(N185),
	.B(N169),
	.C(n2726),
	.D(n2730),
	.OUT(n2729));
   OAI22 U2485 (.OUT(n2731),
	.D(n771),
	.C(n2733),
	.B(n2729),
	.A(n2732));
   AOI22 U2486 (.A(N187),
	.B(N171),
	.C(n2731),
	.D(n2735),
	.OUT(n2734));
   OAI22 U2487 (.OUT(n2736),
	.D(n773),
	.C(n2738),
	.B(n2734),
	.A(n2737));
   AOI22 U2488 (.A(N189),
	.B(N173),
	.C(n2736),
	.D(n2740),
	.OUT(n2739));
   AOI22 U2489 (.A(N190),
	.B(N174),
	.C(n2742),
	.D(n2743),
	.OUT(n2741));
   OAI22 U2490 (.OUT(n2466),
	.D(n776),
	.C(n2106),
	.B(n2741),
	.A(n2105));
   AOI21 U2491 (.OUT(n2744),
	.C(n2234),
	.B(n2109),
	.A(n2112));
   INVERTER U2492 (.IN(n2116),
	.OUT(n2120));
   OAI21 U2493 (.OUT(n2121),
	.C(n2745),
	.B(n2116),
	.A(N215));
   INVERTER U2494 (.IN(n789),
	.OUT(n2123));
   INVERTER U2495 (.IN(n806),
	.OUT(n2468));
   OAI22 U2496 (.OUT(n2467),
	.D(n2221),
	.C(n2137),
	.B(n805),
	.A(n2468));
   OAI21 U2497 (.OUT(n2746),
	.C(n1373),
	.B(n1372),
	.A(n2476));
   OAI21 U2498 (.OUT(n2747),
	.C(n2746),
	.B(n2138),
	.A(n2469));
   OAI21 U2499 (.OUT(n2748),
	.C(n2747),
	.B(N83),
	.A(N99));
   AOI21 U2500 (.OUT(n2749),
	.C(n2750),
	.B(N83),
	.A(N99));
   OAI22 U2501 (.OUT(n2751),
	.D(n807),
	.C(n2753),
	.B(n2749),
	.A(n2752));
   AOI22 U2502 (.A(N101),
	.B(N85),
	.C(n2751),
	.D(n2755),
	.OUT(n2754));
   OAI22 U2503 (.OUT(n2756),
	.D(n809),
	.C(n2758),
	.B(n2754),
	.A(n2757));
   AOI22 U2504 (.A(N103),
	.B(N87),
	.C(n2756),
	.D(n2760),
	.OUT(n2759));
   OAI22 U2505 (.OUT(n2761),
	.D(n811),
	.C(n2763),
	.B(n2759),
	.A(n2762));
   AOI22 U2506 (.A(N105),
	.B(N89),
	.C(n2761),
	.D(n2765),
	.OUT(n2764));
   OAI22 U2507 (.OUT(n2766),
	.D(n813),
	.C(n2768),
	.B(n2764),
	.A(n2767));
   AOI22 U2508 (.A(N107),
	.B(N91),
	.C(n2766),
	.D(n2770),
	.OUT(n2769));
   OAI22 U2509 (.OUT(n2771),
	.D(n815),
	.C(n2773),
	.B(n2769),
	.A(n2772));
   AOI22 U2510 (.A(N109),
	.B(N93),
	.C(n2771),
	.D(n2775),
	.OUT(n2774));
   AOI22 U2511 (.A(N110),
	.B(N94),
	.C(n2777),
	.D(n2778),
	.OUT(n2776));
   OAI22 U2512 (.OUT(n2472),
	.D(n818),
	.C(n2140),
	.B(n2776),
	.A(n2139));
   AOI21 U2513 (.OUT(n2779),
	.C(n2254),
	.B(n2143),
	.A(n2146));
   INVERTER U2514 (.IN(n2150),
	.OUT(n2154));
   OAI21 U2515 (.OUT(n2155),
	.C(n2780),
	.B(n2150),
	.A(N135));
   INVERTER U2516 (.IN(n831),
	.OUT(n2157));
   INVERTER U2517 (.IN(n848),
	.OUT(n2474));
   OAI22 U2518 (.OUT(n2473),
	.D(n2241),
	.C(n2171),
	.B(n847),
	.A(n2474));
   XOR2 U2519 (.A(n859),
	.B(n2259),
	.OUT(n2781));
   XOR2 U2520 (.A(n853),
	.B(n2261),
	.OUT(n865));
   XOR2 U2521 (.A(n849),
	.B(n2263),
	.OUT(n856));
   XOR2 U2522 (.A(n855),
	.B(n2265),
	.OUT(n885));
   XOR2 U2523 (.A(n2782),
	.B(n2478),
	.OUT(n868));
   XOR2 U2524 (.A(n867),
	.B(n2266),
	.OUT(n871));
   XOR2 U2525 (.A(n2783),
	.B(n2480),
	.OUT(n874));
   XOR2 U2526 (.A(n873),
	.B(n2268),
	.OUT(n2499));
   XOR2 U2527 (.A(n862),
	.B(n2269),
	.OUT(n891));
   XOR2 U2528 (.A(n864),
	.B(n2271),
	.OUT(n894));
   XOR2 U2529 (.A(n2784),
	.B(n2273),
	.OUT(n207));
   XOR2 U2530 (.A(n879),
	.B(n2274),
	.OUT(n1442));
   XOR2 U2531 (.A(n881),
	.B(n2276),
	.OUT(n1448));
   XOR2 U2532 (.A(n884),
	.B(n2277),
	.OUT(n209));
   XOR2 U2533 (.A(n2785),
	.B(n2488),
	.OUT(n897));
   XOR2 U2534 (.A(n2786),
	.B(n2490),
	.OUT(n899));
   XOR2 U2535 (.A(n2787),
	.B(n2494),
	.OUT(n198));
   XOR2 U2536 (.A(n896),
	.B(n2278),
	.OUT(n203));
   XOR2 U2537 (.A(n916),
	.B(n2281),
	.OUT(n2788));
   XOR2 U2538 (.A(n910),
	.B(n2283),
	.OUT(n922));
   XOR2 U2539 (.A(n906),
	.B(n2285),
	.OUT(n913));
   XOR2 U2540 (.A(n912),
	.B(n2287),
	.OUT(n942));
   XOR2 U2541 (.A(n2789),
	.B(n2500),
	.OUT(n925));
   XOR2 U2542 (.A(n924),
	.B(n2288),
	.OUT(n928));
   XOR2 U2543 (.A(n2790),
	.B(n2502),
	.OUT(n931));
   XOR2 U2544 (.A(n930),
	.B(n2290),
	.OUT(n2521));
   XOR2 U2545 (.A(n919),
	.B(n2291),
	.OUT(n948));
   XOR2 U2546 (.A(n921),
	.B(n2293),
	.OUT(n951));
   XOR2 U2547 (.A(n2791),
	.B(n2295),
	.OUT(n191));
   XOR2 U2548 (.A(n936),
	.B(n2296),
	.OUT(n1519));
   XOR2 U2549 (.A(n938),
	.B(n2298),
	.OUT(n1525));
   XOR2 U2550 (.A(n941),
	.B(n2299),
	.OUT(n193));
   XOR2 U2551 (.A(n2792),
	.B(n2510),
	.OUT(n954));
   XOR2 U2552 (.A(n2793),
	.B(n2512),
	.OUT(n956));
   XOR2 U2553 (.A(n2794),
	.B(n2516),
	.OUT(n182));
   XOR2 U2554 (.A(n953),
	.B(n2300),
	.OUT(n187));
   XOR2 U2555 (.A(n973),
	.B(n2303),
	.OUT(n2795));
   XOR2 U2556 (.A(n967),
	.B(n2305),
	.OUT(n979));
   XOR2 U2557 (.A(n963),
	.B(n2307),
	.OUT(n970));
   XOR2 U2558 (.A(n969),
	.B(n2309),
	.OUT(n999));
   XOR2 U2559 (.A(n2796),
	.B(n2522),
	.OUT(n982));
   XOR2 U2560 (.A(n981),
	.B(n2310),
	.OUT(n985));
   XOR2 U2561 (.A(n2797),
	.B(n2524),
	.OUT(n988));
   XOR2 U2562 (.A(n987),
	.B(n2312),
	.OUT(n2543));
   XOR2 U2563 (.A(n976),
	.B(n2313),
	.OUT(n1005));
   XOR2 U2564 (.A(n978),
	.B(n2315),
	.OUT(n1008));
   XOR2 U2565 (.A(n2798),
	.B(n2317),
	.OUT(n175));
   XOR2 U2566 (.A(n993),
	.B(n2318),
	.OUT(n1596));
   XOR2 U2567 (.A(n995),
	.B(n2320),
	.OUT(n1602));
   XOR2 U2568 (.A(n998),
	.B(n2321),
	.OUT(n177));
   XOR2 U2569 (.A(n2799),
	.B(n2532),
	.OUT(n1011));
   XOR2 U2570 (.A(n2800),
	.B(n2534),
	.OUT(n1013));
   XOR2 U2571 (.A(n2801),
	.B(n2538),
	.OUT(n166));
   XOR2 U2572 (.A(n1010),
	.B(n2322),
	.OUT(n171));
   XOR2 U2573 (.A(n1030),
	.B(n2325),
	.OUT(n2802));
   XOR2 U2574 (.A(n1024),
	.B(n2327),
	.OUT(n1036));
   XOR2 U2575 (.A(n1020),
	.B(n2329),
	.OUT(n1027));
   XOR2 U2576 (.A(n1026),
	.B(n2331),
	.OUT(n1056));
   XOR2 U2577 (.A(n2803),
	.B(n2544),
	.OUT(n1039));
   XOR2 U2578 (.A(n1038),
	.B(n2332),
	.OUT(n1042));
   XOR2 U2579 (.A(n2804),
	.B(n2546),
	.OUT(n1045));
   XOR2 U2580 (.A(n1044),
	.B(n2334),
	.OUT(n2565));
   XOR2 U2581 (.A(n1033),
	.B(n2335),
	.OUT(n1062));
   XOR2 U2582 (.A(n1035),
	.B(n2337),
	.OUT(n1065));
   XOR2 U2583 (.A(n2805),
	.B(n2339),
	.OUT(n159));
   XOR2 U2584 (.A(n1050),
	.B(n2340),
	.OUT(n1673));
   XOR2 U2585 (.A(n1052),
	.B(n2342),
	.OUT(n1679));
   XOR2 U2586 (.A(n1055),
	.B(n2343),
	.OUT(n161));
   XOR2 U2587 (.A(n2806),
	.B(n2554),
	.OUT(n1068));
   XOR2 U2588 (.A(n2807),
	.B(n2556),
	.OUT(n1070));
   XOR2 U2589 (.A(n2808),
	.B(n2560),
	.OUT(n150));
   XOR2 U2590 (.A(n1067),
	.B(n2344),
	.OUT(n155));
   XOR2 U2591 (.A(n1087),
	.B(n2347),
	.OUT(n2809));
   XOR2 U2592 (.A(n1081),
	.B(n2349),
	.OUT(n1093));
   XOR2 U2593 (.A(n1077),
	.B(n2351),
	.OUT(n1084));
   XOR2 U2594 (.A(n1083),
	.B(n2353),
	.OUT(n1113));
   XOR2 U2595 (.A(n2810),
	.B(n2566),
	.OUT(n1096));
   XOR2 U2596 (.A(n1095),
	.B(n2354),
	.OUT(n1099));
   XOR2 U2597 (.A(n2811),
	.B(n2568),
	.OUT(n1102));
   XOR2 U2598 (.A(n1101),
	.B(n2356),
	.OUT(n2587));
   XOR2 U2599 (.A(n1090),
	.B(n2357),
	.OUT(n1119));
   XOR2 U2600 (.A(n1092),
	.B(n2359),
	.OUT(n1122));
   XOR2 U2601 (.A(n2812),
	.B(n2361),
	.OUT(n143));
   XOR2 U2602 (.A(n1107),
	.B(n2362),
	.OUT(n1750));
   XOR2 U2603 (.A(n1109),
	.B(n2364),
	.OUT(n1756));
   XOR2 U2604 (.A(n1112),
	.B(n2365),
	.OUT(n145));
   XOR2 U2605 (.A(n2813),
	.B(n2576),
	.OUT(n1125));
   XOR2 U2606 (.A(n2814),
	.B(n2578),
	.OUT(n1127));
   XOR2 U2607 (.A(n2815),
	.B(n2582),
	.OUT(n134));
   XOR2 U2608 (.A(n1124),
	.B(n2366),
	.OUT(n139));
   XOR2 U2609 (.A(n1144),
	.B(n2369),
	.OUT(n2816));
   XOR2 U2610 (.A(n1138),
	.B(n2371),
	.OUT(n1150));
   XOR2 U2611 (.A(n1134),
	.B(n2373),
	.OUT(n1141));
   XOR2 U2612 (.A(n1140),
	.B(n2375),
	.OUT(n1170));
   XOR2 U2613 (.A(n2817),
	.B(n2588),
	.OUT(n1153));
   XOR2 U2614 (.A(n1152),
	.B(n2376),
	.OUT(n1156));
   XOR2 U2615 (.A(n2818),
	.B(n2590),
	.OUT(n1159));
   XOR2 U2616 (.A(n1158),
	.B(n2378),
	.OUT(n2609));
   XOR2 U2617 (.A(n1147),
	.B(n2379),
	.OUT(n1176));
   XOR2 U2618 (.A(n1149),
	.B(n2381),
	.OUT(n1179));
   XOR2 U2619 (.A(n2819),
	.B(n2383),
	.OUT(n127));
   XOR2 U2620 (.A(n1164),
	.B(n2384),
	.OUT(n1827));
   XOR2 U2621 (.A(n1166),
	.B(n2386),
	.OUT(n1833));
   XOR2 U2622 (.A(n1169),
	.B(n2387),
	.OUT(n129));
   XOR2 U2623 (.A(n2820),
	.B(n2598),
	.OUT(n1182));
   XOR2 U2624 (.A(n2821),
	.B(n2600),
	.OUT(n1184));
   XOR2 U2625 (.A(n2822),
	.B(n2604),
	.OUT(n118));
   XOR2 U2626 (.A(n1181),
	.B(n2388),
	.OUT(n123));
   XOR2 U2627 (.A(n1201),
	.B(n2391),
	.OUT(n2823));
   XOR2 U2628 (.A(n1195),
	.B(n2393),
	.OUT(n1207));
   XOR2 U2629 (.A(n1191),
	.B(n2395),
	.OUT(n1198));
   XOR2 U2630 (.A(n1197),
	.B(n2397),
	.OUT(n1227));
   XOR2 U2631 (.A(n2824),
	.B(n2610),
	.OUT(n1210));
   XOR2 U2632 (.A(n1209),
	.B(n2398),
	.OUT(n1213));
   XOR2 U2633 (.A(n2825),
	.B(n2612),
	.OUT(n1216));
   XOR2 U2634 (.A(n1215),
	.B(n2400),
	.OUT(n2631));
   XOR2 U2635 (.A(n1204),
	.B(n2401),
	.OUT(n1233));
   XOR2 U2636 (.A(n1206),
	.B(n2403),
	.OUT(n1236));
   XOR2 U2637 (.A(n2826),
	.B(n2405),
	.OUT(n111));
   XOR2 U2638 (.A(n1221),
	.B(n2406),
	.OUT(n1904));
   XOR2 U2639 (.A(n1223),
	.B(n2408),
	.OUT(n1910));
   XOR2 U2640 (.A(n1226),
	.B(n2409),
	.OUT(n113));
   XOR2 U2641 (.A(n2827),
	.B(n2620),
	.OUT(n1239));
   XOR2 U2642 (.A(n2828),
	.B(n2622),
	.OUT(n1241));
   XOR2 U2643 (.A(n2829),
	.B(n2626),
	.OUT(n102));
   XOR2 U2644 (.A(n1238),
	.B(n2410),
	.OUT(n107));
   XOR2 U2645 (.A(n1258),
	.B(n2413),
	.OUT(n2830));
   XOR2 U2646 (.A(n1252),
	.B(n2415),
	.OUT(n1264));
   XOR2 U2647 (.A(n1248),
	.B(n2417),
	.OUT(n1255));
   XOR2 U2648 (.A(n1254),
	.B(n2419),
	.OUT(n1284));
   XOR2 U2649 (.A(n2831),
	.B(n2632),
	.OUT(n1267));
   XOR2 U2650 (.A(n1266),
	.B(n2420),
	.OUT(n1270));
   XOR2 U2651 (.A(n2832),
	.B(n2634),
	.OUT(n1273));
   XOR2 U2652 (.A(n1272),
	.B(n2422),
	.OUT(n2653));
   XOR2 U2653 (.A(n1261),
	.B(n2423),
	.OUT(n1290));
   XOR2 U2654 (.A(n1263),
	.B(n2425),
	.OUT(n1293));
   XOR2 U2655 (.A(n2833),
	.B(n2427),
	.OUT(n95));
   XOR2 U2656 (.A(n1278),
	.B(n2428),
	.OUT(n1981));
   XOR2 U2657 (.A(n1280),
	.B(n2430),
	.OUT(n1987));
   XOR2 U2658 (.A(n1283),
	.B(n2431),
	.OUT(n97));
   XOR2 U2659 (.A(n2834),
	.B(n2642),
	.OUT(n1296));
   XOR2 U2660 (.A(n2835),
	.B(n2644),
	.OUT(n1298));
   XOR2 U2661 (.A(n2836),
	.B(n2648),
	.OUT(n86));
   XOR2 U2662 (.A(n1295),
	.B(n2432),
	.OUT(n91));
   XOR2 U2663 (.A(n1315),
	.B(n2435),
	.OUT(n2837));
   XOR2 U2664 (.A(n1309),
	.B(n2437),
	.OUT(n1321));
   XOR2 U2665 (.A(n1305),
	.B(n2439),
	.OUT(n1312));
   XOR2 U2666 (.A(n1311),
	.B(n2441),
	.OUT(n1341));
   XOR2 U2667 (.A(n2838),
	.B(n2654),
	.OUT(n1324));
   XOR2 U2668 (.A(n1323),
	.B(n2442),
	.OUT(n1327));
   XOR2 U2669 (.A(n2839),
	.B(n2656),
	.OUT(n1330));
   XOR2 U2670 (.A(n1329),
	.B(n2444),
	.OUT(n2675));
   XOR2 U2671 (.A(n1318),
	.B(n2445),
	.OUT(n1347));
   XOR2 U2672 (.A(n1320),
	.B(n2447),
	.OUT(n1350));
   XOR2 U2673 (.A(n2840),
	.B(n2449),
	.OUT(n79));
   XOR2 U2674 (.A(n1335),
	.B(n2450),
	.OUT(n2058));
   XOR2 U2675 (.A(n1337),
	.B(n2452),
	.OUT(n2064));
   XOR2 U2676 (.A(n1340),
	.B(n2453),
	.OUT(n81));
   XOR2 U2677 (.A(n2841),
	.B(n2664),
	.OUT(n1353));
   XOR2 U2678 (.A(n2842),
	.B(n2666),
	.OUT(n1355));
   XOR2 U2679 (.A(n2843),
	.B(n2670),
	.OUT(n70));
   XOR2 U2680 (.A(n1352),
	.B(n2454),
	.OUT(n75));
   INVERTER U2681 (.IN(n1362),
	.OUT(n2457));
   XOR2 U2682 (.A(n2677),
	.B(n2458),
	.OUT(n2077));
   XOR2 U2683 (.A(n2844),
	.B(n2679),
	.OUT(n2214));
   XOR2 U2684 (.A(n2845),
	.B(n2681),
	.OUT(n2081));
   XOR2 U2685 (.A(n2846),
	.B(n2684),
	.OUT(n2084));
   XOR2 U2686 (.A(n2847),
	.B(n2686),
	.OUT(n2710));
   XOR2 U2687 (.A(n2848),
	.B(n2689),
	.OUT(n2090));
   XOR2 U2688 (.A(n2849),
	.B(n2691),
	.OUT(n2092));
   XOR2 U2689 (.A(n2850),
	.B(n2694),
	.OUT(n2094));
   XOR2 U2690 (.A(n2851),
	.B(n2696),
	.OUT(n2096));
   XOR2 U2691 (.A(n2852),
	.B(n2699),
	.OUT(n2098));
   XOR2 U2692 (.A(n2853),
	.B(n2701),
	.OUT(n2100));
   XOR2 U2693 (.A(n2854),
	.B(n2704),
	.OUT(n2102));
   XOR2 U2694 (.A(n2855),
	.B(n2706),
	.OUT(n2201));
   INVERTER U2695 (.IN(n1367),
	.OUT(n2463));
   XOR2 U2696 (.A(n2712),
	.B(n2464),
	.OUT(n2111));
   XOR2 U2697 (.A(n2856),
	.B(n2714),
	.OUT(n2234));
   XOR2 U2698 (.A(n2857),
	.B(n2716),
	.OUT(n2115));
   XOR2 U2699 (.A(n2858),
	.B(n2719),
	.OUT(n2118));
   XOR2 U2700 (.A(n2859),
	.B(n2721),
	.OUT(n2745));
   XOR2 U2701 (.A(n2860),
	.B(n2724),
	.OUT(n2124));
   XOR2 U2702 (.A(n2861),
	.B(n2726),
	.OUT(n2126));
   XOR2 U2703 (.A(n2862),
	.B(n2729),
	.OUT(n2128));
   XOR2 U2704 (.A(n2863),
	.B(n2731),
	.OUT(n2130));
   XOR2 U2705 (.A(n2864),
	.B(n2734),
	.OUT(n2132));
   XOR2 U2706 (.A(n2865),
	.B(n2736),
	.OUT(n2134));
   XOR2 U2707 (.A(n2866),
	.B(n2739),
	.OUT(n2136));
   XOR2 U2708 (.A(n2867),
	.B(n2741),
	.OUT(n2221));
   INVERTER U2709 (.IN(n1372),
	.OUT(n2469));
   XOR2 U2710 (.A(n2747),
	.B(n2470),
	.OUT(n2145));
   XOR2 U2711 (.A(n2868),
	.B(n2749),
	.OUT(n2254));
   XOR2 U2712 (.A(n2869),
	.B(n2751),
	.OUT(n2149));
   XOR2 U2713 (.A(n2870),
	.B(n2754),
	.OUT(n2152));
   XOR2 U2714 (.A(n2871),
	.B(n2756),
	.OUT(n2780));
   XOR2 U2715 (.A(n2872),
	.B(n2759),
	.OUT(n2158));
   XOR2 U2716 (.A(n2873),
	.B(n2761),
	.OUT(n2160));
   XOR2 U2717 (.A(n2874),
	.B(n2764),
	.OUT(n2162));
   XOR2 U2718 (.A(n2875),
	.B(n2766),
	.OUT(n2164));
   XOR2 U2719 (.A(n2876),
	.B(n2769),
	.OUT(n2166));
   XOR2 U2720 (.A(n2877),
	.B(n2771),
	.OUT(n2168));
   XOR2 U2721 (.A(n2878),
	.B(n2774),
	.OUT(n2170));
   XOR2 U2722 (.A(n2879),
	.B(n2776),
	.OUT(n2241));
   XOR2 U2723 (.A(\mult_21_3/ab[2][7] ),
	.B(\mult_21_3/ab[3][6] ),
	.OUT(n2782));
   XOR2 U2724 (.A(\mult_21_3/ab[3][7] ),
	.B(\mult_21_3/ab[4][6] ),
	.OUT(n2783));
   XOR2 U2725 (.A(\mult_21_3/ab[4][7] ),
	.B(n2492),
	.OUT(n2785));
   XOR2 U2726 (.A(\mult_21_3/ab[5][7] ),
	.B(n256),
	.OUT(n2786));
   XOR2 U2727 (.A(\mult_21_3/ab[6][7] ),
	.B(\mult_21_3/ab[7][6] ),
	.OUT(n2787));
   XOR2 U2728 (.A(\mult_21_2/ab[2][7] ),
	.B(\mult_21_2/ab[3][6] ),
	.OUT(n2789));
   XOR2 U2729 (.A(\mult_21_2/ab[3][7] ),
	.B(\mult_21_2/ab[4][6] ),
	.OUT(n2790));
   XOR2 U2730 (.A(\mult_21_2/ab[4][7] ),
	.B(n2514),
	.OUT(n2792));
   XOR2 U2731 (.A(\mult_21_2/ab[5][7] ),
	.B(n313),
	.OUT(n2793));
   XOR2 U2732 (.A(\mult_21_2/ab[6][7] ),
	.B(\mult_21_2/ab[7][6] ),
	.OUT(n2794));
   XOR2 U2733 (.A(\mult_21/ab[2][7] ),
	.B(\mult_21/ab[3][6] ),
	.OUT(n2796));
   XOR2 U2734 (.A(\mult_21/ab[3][7] ),
	.B(\mult_21/ab[4][6] ),
	.OUT(n2797));
   XOR2 U2735 (.A(\mult_21/ab[4][7] ),
	.B(n2536),
	.OUT(n2799));
   XOR2 U2736 (.A(\mult_21/ab[5][7] ),
	.B(n370),
	.OUT(n2800));
   XOR2 U2737 (.A(\mult_21/ab[6][7] ),
	.B(\mult_21/ab[7][6] ),
	.OUT(n2801));
   XOR2 U2738 (.A(\mult_20_3/ab[2][7] ),
	.B(\mult_20_3/ab[3][6] ),
	.OUT(n2803));
   XOR2 U2739 (.A(\mult_20_3/ab[3][7] ),
	.B(\mult_20_3/ab[4][6] ),
	.OUT(n2804));
   XOR2 U2740 (.A(\mult_20_3/ab[4][7] ),
	.B(n2558),
	.OUT(n2806));
   XOR2 U2741 (.A(\mult_20_3/ab[5][7] ),
	.B(n427),
	.OUT(n2807));
   XOR2 U2742 (.A(\mult_20_3/ab[6][7] ),
	.B(\mult_20_3/ab[7][6] ),
	.OUT(n2808));
   XOR2 U2743 (.A(\mult_20_2/ab[2][7] ),
	.B(\mult_20_2/ab[3][6] ),
	.OUT(n2810));
   XOR2 U2744 (.A(\mult_20_2/ab[3][7] ),
	.B(\mult_20_2/ab[4][6] ),
	.OUT(n2811));
   XOR2 U2745 (.A(\mult_20_2/ab[4][7] ),
	.B(n2580),
	.OUT(n2813));
   XOR2 U2746 (.A(\mult_20_2/ab[5][7] ),
	.B(n484),
	.OUT(n2814));
   XOR2 U2747 (.A(\mult_20_2/ab[6][7] ),
	.B(\mult_20_2/ab[7][6] ),
	.OUT(n2815));
   XOR2 U2748 (.A(\mult_20/ab[2][7] ),
	.B(\mult_20/ab[3][6] ),
	.OUT(n2817));
   XOR2 U2749 (.A(\mult_20/ab[3][7] ),
	.B(\mult_20/ab[4][6] ),
	.OUT(n2818));
   XOR2 U2750 (.A(\mult_20/ab[4][7] ),
	.B(n2602),
	.OUT(n2820));
   XOR2 U2751 (.A(\mult_20/ab[5][7] ),
	.B(n541),
	.OUT(n2821));
   XOR2 U2752 (.A(\mult_20/ab[6][7] ),
	.B(\mult_20/ab[7][6] ),
	.OUT(n2822));
   XOR2 U2753 (.A(\mult_19_3/ab[2][7] ),
	.B(\mult_19_3/ab[3][6] ),
	.OUT(n2824));
   XOR2 U2754 (.A(\mult_19_3/ab[3][7] ),
	.B(\mult_19_3/ab[4][6] ),
	.OUT(n2825));
   XOR2 U2755 (.A(\mult_19_3/ab[4][7] ),
	.B(n2624),
	.OUT(n2827));
   XOR2 U2756 (.A(\mult_19_3/ab[5][7] ),
	.B(n598),
	.OUT(n2828));
   XOR2 U2757 (.A(\mult_19_3/ab[6][7] ),
	.B(\mult_19_3/ab[7][6] ),
	.OUT(n2829));
   XOR2 U2758 (.A(\mult_19_2/ab[2][7] ),
	.B(\mult_19_2/ab[3][6] ),
	.OUT(n2831));
   XOR2 U2759 (.A(\mult_19_2/ab[3][7] ),
	.B(\mult_19_2/ab[4][6] ),
	.OUT(n2832));
   XOR2 U2760 (.A(\mult_19_2/ab[4][7] ),
	.B(n2646),
	.OUT(n2834));
   XOR2 U2761 (.A(\mult_19_2/ab[5][7] ),
	.B(n655),
	.OUT(n2835));
   XOR2 U2762 (.A(\mult_19_2/ab[6][7] ),
	.B(\mult_19_2/ab[7][6] ),
	.OUT(n2836));
   XOR2 U2763 (.A(\mult_19/ab[2][7] ),
	.B(\mult_19/ab[3][6] ),
	.OUT(n2838));
   XOR2 U2764 (.A(\mult_19/ab[3][7] ),
	.B(\mult_19/ab[4][6] ),
	.OUT(n2839));
   XOR2 U2765 (.A(\mult_19/ab[4][7] ),
	.B(n2668),
	.OUT(n2841));
   XOR2 U2766 (.A(\mult_19/ab[5][7] ),
	.B(n712),
	.OUT(n2842));
   XOR2 U2767 (.A(\mult_19/ab[6][7] ),
	.B(\mult_19/ab[7][6] ),
	.OUT(n2843));
   XOR2 U2768 (.A(N20),
	.B(N4),
	.OUT(n2844));
   XOR2 U2769 (.A(N21),
	.B(N5),
	.OUT(n2845));
   XOR2 U2770 (.A(N22),
	.B(N6),
	.OUT(n2846));
   XOR2 U2771 (.A(N23),
	.B(N7),
	.OUT(n2847));
   XOR2 U2772 (.A(N24),
	.B(N8),
	.OUT(n2848));
   XOR2 U2773 (.A(N25),
	.B(N9),
	.OUT(n2849));
   XOR2 U2774 (.A(N26),
	.B(N10),
	.OUT(n2850));
   XOR2 U2775 (.A(N27),
	.B(N11),
	.OUT(n2851));
   XOR2 U2776 (.A(N28),
	.B(N12),
	.OUT(n2852));
   XOR2 U2777 (.A(N29),
	.B(N13),
	.OUT(n2853));
   XOR2 U2778 (.A(N30),
	.B(N14),
	.OUT(n2854));
   XOR2 U2779 (.A(N31),
	.B(N15),
	.OUT(n2855));
   XOR2 U2780 (.A(N180),
	.B(N164),
	.OUT(n2856));
   XOR2 U2781 (.A(N181),
	.B(N165),
	.OUT(n2857));
   XOR2 U2782 (.A(N182),
	.B(N166),
	.OUT(n2858));
   XOR2 U2783 (.A(N183),
	.B(N167),
	.OUT(n2859));
   XOR2 U2784 (.A(N184),
	.B(N168),
	.OUT(n2860));
   XOR2 U2785 (.A(N185),
	.B(N169),
	.OUT(n2861));
   XOR2 U2786 (.A(N186),
	.B(N170),
	.OUT(n2862));
   XOR2 U2787 (.A(N187),
	.B(N171),
	.OUT(n2863));
   XOR2 U2788 (.A(N188),
	.B(N172),
	.OUT(n2864));
   XOR2 U2789 (.A(N189),
	.B(N173),
	.OUT(n2865));
   XOR2 U2790 (.A(N190),
	.B(N174),
	.OUT(n2866));
   XOR2 U2791 (.A(N191),
	.B(N175),
	.OUT(n2867));
   XOR2 U2792 (.A(N100),
	.B(N84),
	.OUT(n2868));
   XOR2 U2793 (.A(N101),
	.B(N85),
	.OUT(n2869));
   XOR2 U2794 (.A(N102),
	.B(N86),
	.OUT(n2870));
   XOR2 U2795 (.A(N103),
	.B(N87),
	.OUT(n2871));
   XOR2 U2796 (.A(N104),
	.B(N88),
	.OUT(n2872));
   XOR2 U2797 (.A(N105),
	.B(N89),
	.OUT(n2873));
   XOR2 U2798 (.A(N106),
	.B(N90),
	.OUT(n2874));
   XOR2 U2799 (.A(N107),
	.B(N91),
	.OUT(n2875));
   XOR2 U2800 (.A(N108),
	.B(N92),
	.OUT(n2876));
   XOR2 U2801 (.A(N109),
	.B(N93),
	.OUT(n2877));
   XOR2 U2802 (.A(N110),
	.B(N94),
	.OUT(n2878));
   XOR2 U2803 (.A(N111),
	.B(N95),
	.OUT(n2879));
   INVERTER U2804 (.IN(n1377),
	.OUT(n229));
   INVERTER U2805 (.IN(n230),
	.OUT(n1386));
   INVERTER U2806 (.IN(n1421),
	.OUT(n237));
   INVERTER U2807 (.IN(n1434),
	.OUT(n245));
   INVERTER U2808 (.IN(n250),
	.OUT(n2487));
   INVERTER U2809 (.IN(n884),
	.OUT(n2485));
   INVERTER U2810 (.IN(n252),
	.OUT(n2489));
   INVERTER U2811 (.IN(n2493),
	.OUT(n2494));
   INVERTER U2812 (.IN(n257),
	.OUT(n2495));
   INVERTER U2813 (.IN(n258),
	.OUT(n1450));
   INVERTER U2814 (.IN(n196),
	.OUT(\mult_21_3/A2[12] ));
   INVERTER U2815 (.IN(n199),
	.OUT(\mult_21_3/A2[11] ));
   INVERTER U2816 (.IN(n265),
	.OUT(n2498));
   INVERTER U2817 (.IN(n1454),
	.OUT(n286));
   INVERTER U2818 (.IN(n287),
	.OUT(n1463));
   INVERTER U2819 (.IN(n1498),
	.OUT(n294));
   INVERTER U2820 (.IN(n1511),
	.OUT(n302));
   INVERTER U2821 (.IN(n307),
	.OUT(n2509));
   INVERTER U2822 (.IN(n941),
	.OUT(n2507));
   INVERTER U2823 (.IN(n309),
	.OUT(n2511));
   INVERTER U2824 (.IN(n2515),
	.OUT(n2516));
   INVERTER U2825 (.IN(n314),
	.OUT(n2517));
   INVERTER U2826 (.IN(n315),
	.OUT(n1527));
   INVERTER U2827 (.IN(n180),
	.OUT(\mult_21_2/A2[12] ));
   INVERTER U2828 (.IN(n183),
	.OUT(\mult_21_2/A2[11] ));
   INVERTER U2829 (.IN(n322),
	.OUT(n2520));
   INVERTER U2830 (.IN(n1531),
	.OUT(n343));
   INVERTER U2831 (.IN(n344),
	.OUT(n1540));
   INVERTER U2832 (.IN(n1575),
	.OUT(n351));
   INVERTER U2833 (.IN(n1588),
	.OUT(n359));
   INVERTER U2834 (.IN(n364),
	.OUT(n2531));
   INVERTER U2835 (.IN(n998),
	.OUT(n2529));
   INVERTER U2836 (.IN(n366),
	.OUT(n2533));
   INVERTER U2837 (.IN(n2537),
	.OUT(n2538));
   INVERTER U2838 (.IN(n371),
	.OUT(n2539));
   INVERTER U2839 (.IN(n372),
	.OUT(n1604));
   INVERTER U2840 (.IN(n164),
	.OUT(\mult_21/A2[12] ));
   INVERTER U2841 (.IN(n167),
	.OUT(\mult_21/A2[11] ));
   INVERTER U2842 (.IN(n379),
	.OUT(n2542));
   INVERTER U2843 (.IN(n1608),
	.OUT(n400));
   INVERTER U2844 (.IN(n401),
	.OUT(n1617));
   INVERTER U2845 (.IN(n1652),
	.OUT(n408));
   INVERTER U2846 (.IN(n1665),
	.OUT(n416));
   INVERTER U2847 (.IN(n421),
	.OUT(n2553));
   INVERTER U2848 (.IN(n1055),
	.OUT(n2551));
   INVERTER U2849 (.IN(n423),
	.OUT(n2555));
   INVERTER U2850 (.IN(n2559),
	.OUT(n2560));
   INVERTER U2851 (.IN(n428),
	.OUT(n2561));
   INVERTER U2852 (.IN(n429),
	.OUT(n1681));
   INVERTER U2853 (.IN(n148),
	.OUT(\mult_20_3/A2[12] ));
   INVERTER U2854 (.IN(n151),
	.OUT(\mult_20_3/A2[11] ));
   INVERTER U2855 (.IN(n436),
	.OUT(n2564));
   INVERTER U2856 (.IN(n1685),
	.OUT(n457));
   INVERTER U2857 (.IN(n458),
	.OUT(n1694));
   INVERTER U2858 (.IN(n1729),
	.OUT(n465));
   INVERTER U2859 (.IN(n1742),
	.OUT(n473));
   INVERTER U2860 (.IN(n478),
	.OUT(n2575));
   INVERTER U2861 (.IN(n1112),
	.OUT(n2573));
   INVERTER U2862 (.IN(n480),
	.OUT(n2577));
   INVERTER U2863 (.IN(n2581),
	.OUT(n2582));
   INVERTER U2864 (.IN(n485),
	.OUT(n2583));
   INVERTER U2865 (.IN(n486),
	.OUT(n1758));
   INVERTER U2866 (.IN(n132),
	.OUT(\mult_20_2/A2[12] ));
   INVERTER U2867 (.IN(n135),
	.OUT(\mult_20_2/A2[11] ));
   INVERTER U2868 (.IN(n493),
	.OUT(n2586));
   INVERTER U2869 (.IN(n1762),
	.OUT(n514));
   INVERTER U2870 (.IN(n515),
	.OUT(n1771));
   INVERTER U2871 (.IN(n1806),
	.OUT(n522));
   INVERTER U2872 (.IN(n1819),
	.OUT(n530));
   INVERTER U2873 (.IN(n535),
	.OUT(n2597));
   INVERTER U2874 (.IN(n1169),
	.OUT(n2595));
   INVERTER U2875 (.IN(n537),
	.OUT(n2599));
   INVERTER U2876 (.IN(n2603),
	.OUT(n2604));
   INVERTER U2877 (.IN(n542),
	.OUT(n2605));
   INVERTER U2878 (.IN(n543),
	.OUT(n1835));
   INVERTER U2879 (.IN(n116),
	.OUT(\mult_20/A2[12] ));
   INVERTER U2880 (.IN(n119),
	.OUT(\mult_20/A2[11] ));
   INVERTER U2881 (.IN(n550),
	.OUT(n2608));
   INVERTER U2882 (.IN(n1839),
	.OUT(n571));
   INVERTER U2883 (.IN(n572),
	.OUT(n1848));
   INVERTER U2884 (.IN(n1883),
	.OUT(n579));
   INVERTER U2885 (.IN(n1896),
	.OUT(n587));
   INVERTER U2886 (.IN(n592),
	.OUT(n2619));
   INVERTER U2887 (.IN(n1226),
	.OUT(n2617));
   INVERTER U2888 (.IN(n594),
	.OUT(n2621));
   INVERTER U2889 (.IN(n2625),
	.OUT(n2626));
   INVERTER U2890 (.IN(n599),
	.OUT(n2627));
   INVERTER U2891 (.IN(n600),
	.OUT(n1912));
   INVERTER U2892 (.IN(n100),
	.OUT(\mult_19_3/A2[12] ));
   INVERTER U2893 (.IN(n103),
	.OUT(\mult_19_3/A2[11] ));
   INVERTER U2894 (.IN(n607),
	.OUT(n2630));
   INVERTER U2895 (.IN(n1916),
	.OUT(n628));
   INVERTER U2896 (.IN(n629),
	.OUT(n1925));
   INVERTER U2897 (.IN(n1960),
	.OUT(n636));
   INVERTER U2898 (.IN(n1973),
	.OUT(n644));
   INVERTER U2899 (.IN(n649),
	.OUT(n2641));
   INVERTER U2900 (.IN(n1283),
	.OUT(n2639));
   INVERTER U2901 (.IN(n651),
	.OUT(n2643));
   INVERTER U2902 (.IN(n2647),
	.OUT(n2648));
   INVERTER U2903 (.IN(n656),
	.OUT(n2649));
   INVERTER U2904 (.IN(n657),
	.OUT(n1989));
   INVERTER U2905 (.IN(n84),
	.OUT(\mult_19_2/A2[12] ));
   INVERTER U2906 (.IN(n87),
	.OUT(\mult_19_2/A2[11] ));
   INVERTER U2907 (.IN(n664),
	.OUT(n2652));
   INVERTER U2908 (.IN(n1993),
	.OUT(n685));
   INVERTER U2909 (.IN(n686),
	.OUT(n2002));
   INVERTER U2910 (.IN(n2037),
	.OUT(n693));
   INVERTER U2911 (.IN(n2050),
	.OUT(n701));
   INVERTER U2912 (.IN(n706),
	.OUT(n2663));
   INVERTER U2913 (.IN(n1340),
	.OUT(n2661));
   INVERTER U2914 (.IN(n708),
	.OUT(n2665));
   INVERTER U2915 (.IN(n2669),
	.OUT(n2670));
   INVERTER U2916 (.IN(n713),
	.OUT(n2671));
   INVERTER U2917 (.IN(n714),
	.OUT(n2066));
   INVERTER U2918 (.IN(n68),
	.OUT(\mult_19/A2[12] ));
   INVERTER U2919 (.IN(n71),
	.OUT(\mult_19/A2[11] ));
   INVERTER U2920 (.IN(n721),
	.OUT(n2674));
   INVERTER U2921 (.IN(n2678),
	.OUT(n2680));
   INVERTER U2922 (.IN(n724),
	.OUT(n2685));
   INVERTER U2923 (.IN(n726),
	.OUT(n2690));
   INVERTER U2924 (.IN(n728),
	.OUT(n2695));
   INVERTER U2925 (.IN(n730),
	.OUT(n2700));
   INVERTER U2926 (.IN(n732),
	.OUT(n2705));
   INVERTER U2927 (.IN(n2704),
	.OUT(n2707));
   INVERTER U2928 (.IN(n733),
	.OUT(n2708));
   INVERTER U2929 (.IN(n2073),
	.OUT(n736));
   INVERTER U2930 (.IN(n2713),
	.OUT(n2715));
   INVERTER U2931 (.IN(n766),
	.OUT(n2720));
   INVERTER U2932 (.IN(n768),
	.OUT(n2725));
   INVERTER U2933 (.IN(n770),
	.OUT(n2730));
   INVERTER U2934 (.IN(n772),
	.OUT(n2735));
   INVERTER U2935 (.IN(n774),
	.OUT(n2740));
   INVERTER U2936 (.IN(n2739),
	.OUT(n2742));
   INVERTER U2937 (.IN(n775),
	.OUT(n2743));
   INVERTER U2938 (.IN(n2107),
	.OUT(n778));
   INVERTER U2939 (.IN(n2748),
	.OUT(n2750));
   INVERTER U2940 (.IN(n808),
	.OUT(n2755));
   INVERTER U2941 (.IN(n810),
	.OUT(n2760));
   INVERTER U2942 (.IN(n812),
	.OUT(n2765));
   INVERTER U2943 (.IN(n814),
	.OUT(n2770));
   INVERTER U2944 (.IN(n816),
	.OUT(n2775));
   INVERTER U2945 (.IN(n2774),
	.OUT(n2777));
   INVERTER U2946 (.IN(n817),
	.OUT(n2778));
   INVERTER U2947 (.IN(n2141),
	.OUT(n820));
   INVERTER U2948 (.IN(n233),
	.OUT(n1405));
   INVERTER U2949 (.IN(\mult_21_3/ab[6][2] ),
	.OUT(n1406));
   INVERTER U2950 (.IN(n234),
	.OUT(n2483));
   INVERTER U2951 (.IN(n214),
	.OUT(n1416));
   INVERTER U2952 (.IN(n241),
	.OUT(n1432));
   INVERTER U2953 (.IN(\mult_21_3/ab[6][1] ),
	.OUT(n1433));
   INVERTER U2954 (.IN(n242),
	.OUT(n2484));
   INVERTER U2955 (.IN(\mult_21_3/ab[4][7] ),
	.OUT(n2491));
   INVERTER U2956 (.IN(\mult_21_3/ab[5][6] ),
	.OUT(n2492));
   INVERTER U2957 (.IN(n890),
	.OUT(n2486));
   INVERTER U2958 (.IN(n290),
	.OUT(n1482));
   INVERTER U2959 (.IN(\mult_21_2/ab[6][2] ),
	.OUT(n1483));
   INVERTER U2960 (.IN(n291),
	.OUT(n2505));
   INVERTER U2961 (.IN(n271),
	.OUT(n1493));
   INVERTER U2962 (.IN(n298),
	.OUT(n1509));
   INVERTER U2963 (.IN(\mult_21_2/ab[6][1] ),
	.OUT(n1510));
   INVERTER U2964 (.IN(n299),
	.OUT(n2506));
   INVERTER U2965 (.IN(\mult_21_2/ab[4][7] ),
	.OUT(n2513));
   INVERTER U2966 (.IN(\mult_21_2/ab[5][6] ),
	.OUT(n2514));
   INVERTER U2967 (.IN(n947),
	.OUT(n2508));
   INVERTER U2968 (.IN(n347),
	.OUT(n1559));
   INVERTER U2969 (.IN(\mult_21/ab[6][2] ),
	.OUT(n1560));
   INVERTER U2970 (.IN(n348),
	.OUT(n2527));
   INVERTER U2971 (.IN(n328),
	.OUT(n1570));
   INVERTER U2972 (.IN(n355),
	.OUT(n1586));
   INVERTER U2973 (.IN(\mult_21/ab[6][1] ),
	.OUT(n1587));
   INVERTER U2974 (.IN(n356),
	.OUT(n2528));
   INVERTER U2975 (.IN(\mult_21/ab[4][7] ),
	.OUT(n2535));
   INVERTER U2976 (.IN(\mult_21/ab[5][6] ),
	.OUT(n2536));
   INVERTER U2977 (.IN(n1004),
	.OUT(n2530));
   INVERTER U2978 (.IN(n404),
	.OUT(n1636));
   INVERTER U2979 (.IN(\mult_20_3/ab[6][2] ),
	.OUT(n1637));
   INVERTER U2980 (.IN(n405),
	.OUT(n2549));
   INVERTER U2981 (.IN(n385),
	.OUT(n1647));
   INVERTER U2982 (.IN(n412),
	.OUT(n1663));
   INVERTER U2983 (.IN(\mult_20_3/ab[6][1] ),
	.OUT(n1664));
   INVERTER U2984 (.IN(n413),
	.OUT(n2550));
   INVERTER U2985 (.IN(\mult_20_3/ab[4][7] ),
	.OUT(n2557));
   INVERTER U2986 (.IN(\mult_20_3/ab[5][6] ),
	.OUT(n2558));
   INVERTER U2987 (.IN(n1061),
	.OUT(n2552));
   INVERTER U2988 (.IN(n461),
	.OUT(n1713));
   INVERTER U2989 (.IN(\mult_20_2/ab[6][2] ),
	.OUT(n1714));
   INVERTER U2990 (.IN(n462),
	.OUT(n2571));
   INVERTER U2991 (.IN(n442),
	.OUT(n1724));
   INVERTER U2992 (.IN(n469),
	.OUT(n1740));
   INVERTER U2993 (.IN(\mult_20_2/ab[6][1] ),
	.OUT(n1741));
   INVERTER U2994 (.IN(n470),
	.OUT(n2572));
   INVERTER U2995 (.IN(\mult_20_2/ab[4][7] ),
	.OUT(n2579));
   INVERTER U2996 (.IN(\mult_20_2/ab[5][6] ),
	.OUT(n2580));
   INVERTER U2997 (.IN(n1118),
	.OUT(n2574));
   INVERTER U2998 (.IN(n518),
	.OUT(n1790));
   INVERTER U2999 (.IN(\mult_20/ab[6][2] ),
	.OUT(n1791));
   INVERTER U3000 (.IN(n519),
	.OUT(n2593));
   INVERTER U3001 (.IN(n499),
	.OUT(n1801));
   INVERTER U3002 (.IN(n526),
	.OUT(n1817));
   INVERTER U3003 (.IN(\mult_20/ab[6][1] ),
	.OUT(n1818));
   INVERTER U3004 (.IN(n527),
	.OUT(n2594));
   INVERTER U3005 (.IN(\mult_20/ab[4][7] ),
	.OUT(n2601));
   INVERTER U3006 (.IN(\mult_20/ab[5][6] ),
	.OUT(n2602));
   INVERTER U3007 (.IN(n1175),
	.OUT(n2596));
   INVERTER U3008 (.IN(n575),
	.OUT(n1867));
   INVERTER U3009 (.IN(\mult_19_3/ab[6][2] ),
	.OUT(n1868));
   INVERTER U3010 (.IN(n576),
	.OUT(n2615));
   INVERTER U3011 (.IN(n556),
	.OUT(n1878));
   INVERTER U3012 (.IN(n583),
	.OUT(n1894));
   INVERTER U3013 (.IN(\mult_19_3/ab[6][1] ),
	.OUT(n1895));
   INVERTER U3014 (.IN(n584),
	.OUT(n2616));
   INVERTER U3015 (.IN(\mult_19_3/ab[4][7] ),
	.OUT(n2623));
   INVERTER U3016 (.IN(\mult_19_3/ab[5][6] ),
	.OUT(n2624));
   INVERTER U3017 (.IN(n1232),
	.OUT(n2618));
   INVERTER U3018 (.IN(n632),
	.OUT(n1944));
   INVERTER U3019 (.IN(\mult_19_2/ab[6][2] ),
	.OUT(n1945));
   INVERTER U3020 (.IN(n633),
	.OUT(n2637));
   INVERTER U3021 (.IN(n613),
	.OUT(n1955));
   INVERTER U3022 (.IN(n640),
	.OUT(n1971));
   INVERTER U3023 (.IN(\mult_19_2/ab[6][1] ),
	.OUT(n1972));
   INVERTER U3024 (.IN(n641),
	.OUT(n2638));
   INVERTER U3025 (.IN(\mult_19_2/ab[4][7] ),
	.OUT(n2645));
   INVERTER U3026 (.IN(\mult_19_2/ab[5][6] ),
	.OUT(n2646));
   INVERTER U3027 (.IN(n1289),
	.OUT(n2640));
   INVERTER U3028 (.IN(n689),
	.OUT(n2021));
   INVERTER U3029 (.IN(\mult_19/ab[6][2] ),
	.OUT(n2022));
   INVERTER U3030 (.IN(n690),
	.OUT(n2659));
   INVERTER U3031 (.IN(n670),
	.OUT(n2032));
   INVERTER U3032 (.IN(n697),
	.OUT(n2048));
   INVERTER U3033 (.IN(\mult_19/ab[6][1] ),
	.OUT(n2049));
   INVERTER U3034 (.IN(n698),
	.OUT(n2660));
   INVERTER U3035 (.IN(\mult_19/ab[4][7] ),
	.OUT(n2667));
   INVERTER U3036 (.IN(\mult_19/ab[5][6] ),
	.OUT(n2668));
   INVERTER U3037 (.IN(n1346),
	.OUT(n2662));
   INVERTER U3038 (.IN(N20),
	.OUT(n2682));
   INVERTER U3039 (.IN(N4),
	.OUT(n2683));
   INVERTER U3040 (.IN(N22),
	.OUT(n2687));
   INVERTER U3041 (.IN(N6),
	.OUT(n2688));
   INVERTER U3042 (.IN(N24),
	.OUT(n2692));
   INVERTER U3043 (.IN(N8),
	.OUT(n2693));
   INVERTER U3044 (.IN(N26),
	.OUT(n2697));
   INVERTER U3045 (.IN(N10),
	.OUT(n2698));
   INVERTER U3046 (.IN(N28),
	.OUT(n2702));
   INVERTER U3047 (.IN(N12),
	.OUT(n2703));
   INVERTER U3048 (.IN(n740),
	.OUT(n2076));
   INVERTER U3049 (.IN(n741),
	.OUT(n2080));
   INVERTER U3050 (.IN(n748),
	.OUT(n2091));
   INVERTER U3051 (.IN(n753),
	.OUT(n2095));
   INVERTER U3052 (.IN(n758),
	.OUT(n2099));
   INVERTER U3053 (.IN(N180),
	.OUT(n2717));
   INVERTER U3054 (.IN(N164),
	.OUT(n2718));
   INVERTER U3055 (.IN(N182),
	.OUT(n2722));
   INVERTER U3056 (.IN(N166),
	.OUT(n2723));
   INVERTER U3057 (.IN(N184),
	.OUT(n2727));
   INVERTER U3058 (.IN(N168),
	.OUT(n2728));
   INVERTER U3059 (.IN(N186),
	.OUT(n2732));
   INVERTER U3060 (.IN(N170),
	.OUT(n2733));
   INVERTER U3061 (.IN(N188),
	.OUT(n2737));
   INVERTER U3062 (.IN(N172),
	.OUT(n2738));
   INVERTER U3063 (.IN(n782),
	.OUT(n2110));
   INVERTER U3064 (.IN(n783),
	.OUT(n2114));
   INVERTER U3065 (.IN(n790),
	.OUT(n2125));
   INVERTER U3066 (.IN(n795),
	.OUT(n2129));
   INVERTER U3067 (.IN(n800),
	.OUT(n2133));
   INVERTER U3068 (.IN(N100),
	.OUT(n2752));
   INVERTER U3069 (.IN(N84),
	.OUT(n2753));
   INVERTER U3070 (.IN(N102),
	.OUT(n2757));
   INVERTER U3071 (.IN(N86),
	.OUT(n2758));
   INVERTER U3072 (.IN(N104),
	.OUT(n2762));
   INVERTER U3073 (.IN(N88),
	.OUT(n2763));
   INVERTER U3074 (.IN(N106),
	.OUT(n2767));
   INVERTER U3075 (.IN(N90),
	.OUT(n2768));
   INVERTER U3076 (.IN(N108),
	.OUT(n2772));
   INVERTER U3077 (.IN(N92),
	.OUT(n2773));
   INVERTER U3078 (.IN(n824),
	.OUT(n2144));
   INVERTER U3079 (.IN(n825),
	.OUT(n2148));
   INVERTER U3080 (.IN(n832),
	.OUT(n2159));
   INVERTER U3081 (.IN(n837),
	.OUT(n2163));
   INVERTER U3082 (.IN(n842),
	.OUT(n2167));
   INVERTER U3083 (.IN(\mult_21_3/ab[3][6] ),
	.OUT(n2481));
   INVERTER U3084 (.IN(\mult_21_3/ab[2][7] ),
	.OUT(n2482));
   INVERTER U3085 (.IN(\mult_21_2/ab[3][6] ),
	.OUT(n2503));
   INVERTER U3086 (.IN(\mult_21_2/ab[2][7] ),
	.OUT(n2504));
   INVERTER U3087 (.IN(\mult_21/ab[3][6] ),
	.OUT(n2525));
   INVERTER U3088 (.IN(\mult_21/ab[2][7] ),
	.OUT(n2526));
   INVERTER U3089 (.IN(\mult_20_3/ab[3][6] ),
	.OUT(n2547));
   INVERTER U3090 (.IN(\mult_20_3/ab[2][7] ),
	.OUT(n2548));
   INVERTER U3091 (.IN(\mult_20_2/ab[3][6] ),
	.OUT(n2569));
   INVERTER U3092 (.IN(\mult_20_2/ab[2][7] ),
	.OUT(n2570));
   INVERTER U3093 (.IN(\mult_20/ab[3][6] ),
	.OUT(n2591));
   INVERTER U3094 (.IN(\mult_20/ab[2][7] ),
	.OUT(n2592));
   INVERTER U3095 (.IN(\mult_19_3/ab[3][6] ),
	.OUT(n2613));
   INVERTER U3096 (.IN(\mult_19_3/ab[2][7] ),
	.OUT(n2614));
   INVERTER U3097 (.IN(\mult_19_2/ab[3][6] ),
	.OUT(n2635));
   INVERTER U3098 (.IN(\mult_19_2/ab[2][7] ),
	.OUT(n2636));
   INVERTER U3099 (.IN(\mult_19/ab[3][6] ),
	.OUT(n2657));
   INVERTER U3100 (.IN(\mult_19/ab[2][7] ),
	.OUT(n2658));
   INVERTER U3101 (.IN(n2709),
	.OUT(n2079));
   INVERTER U3102 (.IN(n2744),
	.OUT(n2113));
   INVERTER U3103 (.IN(n2779),
	.OUT(n2147));
   INVERTER U3104 (.IN(n239),
	.OUT(n1427));
   INVERTER U3105 (.IN(\mult_21_3/ab[4][1] ),
	.OUT(n1428));
   INVERTER U3106 (.IN(\mult_21_3/ab[5][7] ),
	.OUT(n255));
   INVERTER U3107 (.IN(n296),
	.OUT(n1504));
   INVERTER U3108 (.IN(\mult_21_2/ab[4][1] ),
	.OUT(n1505));
   INVERTER U3109 (.IN(\mult_21_2/ab[5][7] ),
	.OUT(n312));
   INVERTER U3110 (.IN(n353),
	.OUT(n1581));
   INVERTER U3111 (.IN(\mult_21/ab[4][1] ),
	.OUT(n1582));
   INVERTER U3112 (.IN(\mult_21/ab[5][7] ),
	.OUT(n369));
   INVERTER U3113 (.IN(n410),
	.OUT(n1658));
   INVERTER U3114 (.IN(\mult_20_3/ab[4][1] ),
	.OUT(n1659));
   INVERTER U3115 (.IN(\mult_20_3/ab[5][7] ),
	.OUT(n426));
   INVERTER U3116 (.IN(n467),
	.OUT(n1735));
   INVERTER U3117 (.IN(\mult_20_2/ab[4][1] ),
	.OUT(n1736));
   INVERTER U3118 (.IN(\mult_20_2/ab[5][7] ),
	.OUT(n483));
   INVERTER U3119 (.IN(n524),
	.OUT(n1812));
   INVERTER U3120 (.IN(\mult_20/ab[4][1] ),
	.OUT(n1813));
   INVERTER U3121 (.IN(\mult_20/ab[5][7] ),
	.OUT(n540));
   INVERTER U3122 (.IN(n581),
	.OUT(n1889));
   INVERTER U3123 (.IN(\mult_19_3/ab[4][1] ),
	.OUT(n1890));
   INVERTER U3124 (.IN(\mult_19_3/ab[5][7] ),
	.OUT(n597));
   INVERTER U3125 (.IN(n638),
	.OUT(n1966));
   INVERTER U3126 (.IN(\mult_19_2/ab[4][1] ),
	.OUT(n1967));
   INVERTER U3127 (.IN(\mult_19_2/ab[5][7] ),
	.OUT(n654));
   INVERTER U3128 (.IN(n695),
	.OUT(n2043));
   INVERTER U3129 (.IN(\mult_19/ab[4][1] ),
	.OUT(n2044));
   INVERTER U3130 (.IN(\mult_19/ab[5][7] ),
	.OUT(n711));
   INVERTER U3131 (.IN(n228),
	.OUT(n1379));
   INVERTER U3132 (.IN(\mult_21_3/ab[2][3] ),
	.OUT(n222));
   INVERTER U3133 (.IN(n2781),
	.OUT(n882));
   INVERTER U3134 (.IN(\mult_21_3/ab[2][4] ),
	.OUT(n217));
   INVERTER U3135 (.IN(\mult_21_3/ab[2][5] ),
	.OUT(n212));
   INVERTER U3136 (.IN(n2499),
	.OUT(n876));
   INVERTER U3137 (.IN(n236),
	.OUT(n1423));
   INVERTER U3138 (.IN(n870),
	.OUT(n2784));
   INVERTER U3139 (.IN(n244),
	.OUT(n1436));
   INVERTER U3140 (.IN(n893),
	.OUT(n901));
   INVERTER U3141 (.IN(\mult_21_3/ab[6][6] ),
	.OUT(n256));
   INVERTER U3142 (.IN(n260),
	.OUT(n2496));
   INVERTER U3143 (.IN(n904),
	.OUT(\mult_21_3/A1[1] ));
   INVERTER U3144 (.IN(n285),
	.OUT(n1456));
   INVERTER U3145 (.IN(\mult_21_2/ab[2][3] ),
	.OUT(n279));
   INVERTER U3146 (.IN(n2788),
	.OUT(n939));
   INVERTER U3147 (.IN(\mult_21_2/ab[2][4] ),
	.OUT(n274));
   INVERTER U3148 (.IN(\mult_21_2/ab[2][5] ),
	.OUT(n269));
   INVERTER U3149 (.IN(n2521),
	.OUT(n933));
   INVERTER U3150 (.IN(n293),
	.OUT(n1500));
   INVERTER U3151 (.IN(n927),
	.OUT(n2791));
   INVERTER U3152 (.IN(n301),
	.OUT(n1513));
   INVERTER U3153 (.IN(n950),
	.OUT(n958));
   INVERTER U3154 (.IN(\mult_21_2/ab[6][6] ),
	.OUT(n313));
   INVERTER U3155 (.IN(n317),
	.OUT(n2518));
   INVERTER U3156 (.IN(n961),
	.OUT(\mult_21_2/A1[1] ));
   INVERTER U3157 (.IN(n342),
	.OUT(n1533));
   INVERTER U3158 (.IN(\mult_21/ab[2][3] ),
	.OUT(n336));
   INVERTER U3159 (.IN(n2795),
	.OUT(n996));
   INVERTER U3160 (.IN(\mult_21/ab[2][4] ),
	.OUT(n331));
   INVERTER U3161 (.IN(\mult_21/ab[2][5] ),
	.OUT(n326));
   INVERTER U3162 (.IN(n2543),
	.OUT(n990));
   INVERTER U3163 (.IN(n350),
	.OUT(n1577));
   INVERTER U3164 (.IN(n984),
	.OUT(n2798));
   INVERTER U3165 (.IN(n358),
	.OUT(n1590));
   INVERTER U3166 (.IN(n1007),
	.OUT(n1015));
   INVERTER U3167 (.IN(\mult_21/ab[6][6] ),
	.OUT(n370));
   INVERTER U3168 (.IN(n374),
	.OUT(n2540));
   INVERTER U3169 (.IN(n1018),
	.OUT(\mult_21/A1[1] ));
   INVERTER U3170 (.IN(n399),
	.OUT(n1610));
   INVERTER U3171 (.IN(\mult_20_3/ab[2][3] ),
	.OUT(n393));
   INVERTER U3172 (.IN(n2802),
	.OUT(n1053));
   INVERTER U3173 (.IN(\mult_20_3/ab[2][4] ),
	.OUT(n388));
   INVERTER U3174 (.IN(\mult_20_3/ab[2][5] ),
	.OUT(n383));
   INVERTER U3175 (.IN(n2565),
	.OUT(n1047));
   INVERTER U3176 (.IN(n407),
	.OUT(n1654));
   INVERTER U3177 (.IN(n1041),
	.OUT(n2805));
   INVERTER U3178 (.IN(n415),
	.OUT(n1667));
   INVERTER U3179 (.IN(n1064),
	.OUT(n1072));
   INVERTER U3180 (.IN(\mult_20_3/ab[6][6] ),
	.OUT(n427));
   INVERTER U3181 (.IN(n431),
	.OUT(n2562));
   INVERTER U3182 (.IN(n1075),
	.OUT(\mult_20_3/A1[1] ));
   INVERTER U3183 (.IN(n456),
	.OUT(n1687));
   INVERTER U3184 (.IN(\mult_20_2/ab[2][3] ),
	.OUT(n450));
   INVERTER U3185 (.IN(n2809),
	.OUT(n1110));
   INVERTER U3186 (.IN(\mult_20_2/ab[2][4] ),
	.OUT(n445));
   INVERTER U3187 (.IN(\mult_20_2/ab[2][5] ),
	.OUT(n440));
   INVERTER U3188 (.IN(n2587),
	.OUT(n1104));
   INVERTER U3189 (.IN(n464),
	.OUT(n1731));
   INVERTER U3190 (.IN(n1098),
	.OUT(n2812));
   INVERTER U3191 (.IN(n472),
	.OUT(n1744));
   INVERTER U3192 (.IN(n1121),
	.OUT(n1129));
   INVERTER U3193 (.IN(\mult_20_2/ab[6][6] ),
	.OUT(n484));
   INVERTER U3194 (.IN(n488),
	.OUT(n2584));
   INVERTER U3195 (.IN(n1132),
	.OUT(\mult_20_2/A1[1] ));
   INVERTER U3196 (.IN(n513),
	.OUT(n1764));
   INVERTER U3197 (.IN(\mult_20/ab[2][3] ),
	.OUT(n507));
   INVERTER U3198 (.IN(n2816),
	.OUT(n1167));
   INVERTER U3199 (.IN(\mult_20/ab[2][4] ),
	.OUT(n502));
   INVERTER U3200 (.IN(\mult_20/ab[2][5] ),
	.OUT(n497));
   INVERTER U3201 (.IN(n2609),
	.OUT(n1161));
   INVERTER U3202 (.IN(n521),
	.OUT(n1808));
   INVERTER U3203 (.IN(n1155),
	.OUT(n2819));
   INVERTER U3204 (.IN(n529),
	.OUT(n1821));
   INVERTER U3205 (.IN(n1178),
	.OUT(n1186));
   INVERTER U3206 (.IN(\mult_20/ab[6][6] ),
	.OUT(n541));
   INVERTER U3207 (.IN(n545),
	.OUT(n2606));
   INVERTER U3208 (.IN(n1189),
	.OUT(\mult_20/A1[1] ));
   INVERTER U3209 (.IN(n570),
	.OUT(n1841));
   INVERTER U3210 (.IN(\mult_19_3/ab[2][3] ),
	.OUT(n564));
   INVERTER U3211 (.IN(n2823),
	.OUT(n1224));
   INVERTER U3212 (.IN(\mult_19_3/ab[2][4] ),
	.OUT(n559));
   INVERTER U3213 (.IN(\mult_19_3/ab[2][5] ),
	.OUT(n554));
   INVERTER U3214 (.IN(n2631),
	.OUT(n1218));
   INVERTER U3215 (.IN(n578),
	.OUT(n1885));
   INVERTER U3216 (.IN(n1212),
	.OUT(n2826));
   INVERTER U3217 (.IN(n586),
	.OUT(n1898));
   INVERTER U3218 (.IN(n1235),
	.OUT(n1243));
   INVERTER U3219 (.IN(\mult_19_3/ab[6][6] ),
	.OUT(n598));
   INVERTER U3220 (.IN(n602),
	.OUT(n2628));
   INVERTER U3221 (.IN(n1246),
	.OUT(\mult_19_3/A1[1] ));
   INVERTER U3222 (.IN(n627),
	.OUT(n1918));
   INVERTER U3223 (.IN(\mult_19_2/ab[2][3] ),
	.OUT(n621));
   INVERTER U3224 (.IN(n2830),
	.OUT(n1281));
   INVERTER U3225 (.IN(\mult_19_2/ab[2][4] ),
	.OUT(n616));
   INVERTER U3226 (.IN(\mult_19_2/ab[2][5] ),
	.OUT(n611));
   INVERTER U3227 (.IN(n2653),
	.OUT(n1275));
   INVERTER U3228 (.IN(n635),
	.OUT(n1962));
   INVERTER U3229 (.IN(n1269),
	.OUT(n2833));
   INVERTER U3230 (.IN(n643),
	.OUT(n1975));
   INVERTER U3231 (.IN(n1292),
	.OUT(n1300));
   INVERTER U3232 (.IN(\mult_19_2/ab[6][6] ),
	.OUT(n655));
   INVERTER U3233 (.IN(n659),
	.OUT(n2650));
   INVERTER U3234 (.IN(n1303),
	.OUT(\mult_19_2/A1[1] ));
   INVERTER U3235 (.IN(n684),
	.OUT(n1995));
   INVERTER U3236 (.IN(\mult_19/ab[2][3] ),
	.OUT(n678));
   INVERTER U3237 (.IN(n2837),
	.OUT(n1338));
   INVERTER U3238 (.IN(\mult_19/ab[2][4] ),
	.OUT(n673));
   INVERTER U3239 (.IN(\mult_19/ab[2][5] ),
	.OUT(n668));
   INVERTER U3240 (.IN(n2675),
	.OUT(n1332));
   INVERTER U3241 (.IN(n692),
	.OUT(n2039));
   INVERTER U3242 (.IN(n1326),
	.OUT(n2840));
   INVERTER U3243 (.IN(n700),
	.OUT(n2052));
   INVERTER U3244 (.IN(n1349),
	.OUT(n1357));
   INVERTER U3245 (.IN(\mult_19/ab[6][6] ),
	.OUT(n712));
   INVERTER U3246 (.IN(n716),
	.OUT(n2672));
   INVERTER U3247 (.IN(n1360),
	.OUT(\mult_19/A1[1] ));
   INVERTER U3248 (.IN(n735),
	.OUT(n2074));
   INVERTER U3249 (.IN(N51),
	.OUT(n739));
   INVERTER U3250 (.IN(n743),
	.OUT(n2083));
   INVERTER U3251 (.IN(n750),
	.OUT(n2093));
   INVERTER U3252 (.IN(n755),
	.OUT(n2097));
   INVERTER U3253 (.IN(n760),
	.OUT(n2101));
   INVERTER U3254 (.IN(n2710),
	.OUT(n2210));
   INVERTER U3255 (.IN(n2077),
	.OUT(n2216));
   INVERTER U3256 (.IN(n777),
	.OUT(n2108));
   INVERTER U3257 (.IN(N211),
	.OUT(n781));
   INVERTER U3258 (.IN(n785),
	.OUT(n2117));
   INVERTER U3259 (.IN(n792),
	.OUT(n2127));
   INVERTER U3260 (.IN(n797),
	.OUT(n2131));
   INVERTER U3261 (.IN(n802),
	.OUT(n2135));
   INVERTER U3262 (.IN(n2745),
	.OUT(n2230));
   INVERTER U3263 (.IN(n2111),
	.OUT(n2236));
   INVERTER U3264 (.IN(n819),
	.OUT(n2142));
   INVERTER U3265 (.IN(N131),
	.OUT(n823));
   INVERTER U3266 (.IN(n827),
	.OUT(n2151));
   INVERTER U3267 (.IN(n834),
	.OUT(n2161));
   INVERTER U3268 (.IN(n839),
	.OUT(n2165));
   INVERTER U3269 (.IN(n844),
	.OUT(n2169));
   INVERTER U3270 (.IN(n2780),
	.OUT(n2250));
   INVERTER U3271 (.IN(n2145),
	.OUT(n2256));
   INVERTER U3272 (.IN(\mult_19/A1[0] ),
	.OUT(n2880));
   INVERTER U3273 (.IN(n2881),
	.OUT(N3));
   INVERTER U3274 (.IN(\mult_19/A1[1] ),
	.OUT(n2882));
   INVERTER U3275 (.IN(n2883),
	.OUT(N4));
   INVERTER U3276 (.IN(\mult_19/A1[2] ),
	.OUT(n2884));
   INVERTER U3277 (.IN(n2885),
	.OUT(N5));
   INVERTER U3278 (.IN(\mult_19/A1[3] ),
	.OUT(n2886));
   INVERTER U3279 (.IN(n2887),
	.OUT(N6));
   INVERTER U3280 (.IN(\mult_19/A1[4] ),
	.OUT(n2888));
   INVERTER U3281 (.IN(n2889),
	.OUT(N7));
   INVERTER U3282 (.IN(\mult_19/A1[5] ),
	.OUT(n2890));
   INVERTER U3283 (.IN(n2891),
	.OUT(N8));
   INVERTER U3284 (.IN(\mult_19/A1[6] ),
	.OUT(n2892));
   INVERTER U3285 (.IN(n2893),
	.OUT(N9));
   INVERTER U3286 (.IN(\mult_19/A1[7] ),
	.OUT(n2894));
   INVERTER U3287 (.IN(\mult_19/A2[7] ),
	.OUT(n2895));
   INVERTER U3288 (.IN(n2896),
	.OUT(N10));
   INVERTER U3289 (.IN(\mult_19/A1[8] ),
	.OUT(n2897));
   INVERTER U3290 (.IN(\mult_19/A2[8] ),
	.OUT(n2898));
   INVERTER U3291 (.IN(n2899),
	.OUT(\mult_19/FS_1/PG_int[0][2][0] ));
   INVERTER U3292 (.IN(\mult_19/A1[9] ),
	.OUT(n2900));
   INVERTER U3293 (.IN(\mult_19/A2[9] ),
	.OUT(n2901));
   INVERTER U3294 (.IN(n2902),
	.OUT(\mult_19/FS_1/PG_int[0][2][1] ));
   INVERTER U3295 (.IN(n2903),
	.OUT(\mult_19/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3296 (.IN(\mult_19/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2904));
   INVERTER U3297 (.IN(\mult_19/A1[10] ),
	.OUT(n2905));
   INVERTER U3298 (.IN(\mult_19/A2[10] ),
	.OUT(n2906));
   INVERTER U3299 (.IN(n2907),
	.OUT(\mult_19/FS_1/PG_int[0][2][2] ));
   INVERTER U3300 (.IN(n2908),
	.OUT(\mult_19/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3301 (.IN(\mult_19/FS_1/TEMP_G[0][2][1] ),
	.OUT(n2909));
   INVERTER U3302 (.IN(\mult_19/FS_1/C[1][2][1] ),
	.OUT(n2910));
   INVERTER U3303 (.IN(\mult_19/FS_1/P[0][2][1] ),
	.OUT(n2911));
   INVERTER U3304 (.IN(\mult_19/A1[11] ),
	.OUT(n2912));
   INVERTER U3305 (.IN(\mult_19/A2[11] ),
	.OUT(n2913));
   INVERTER U3306 (.IN(n2914),
	.OUT(\mult_19/FS_1/PG_int[0][2][3] ));
   INVERTER U3307 (.IN(\mult_19/FS_1/TEMP_G[0][2][2] ),
	.OUT(n2915));
   INVERTER U3308 (.IN(\mult_19/FS_1/P[0][2][3] ),
	.OUT(n2916));
   INVERTER U3309 (.IN(\mult_19/FS_1/C[1][2][2] ),
	.OUT(n2917));
   INVERTER U3310 (.IN(\mult_19/FS_1/P[0][2][2] ),
	.OUT(n2918));
   INVERTER U3311 (.IN(\mult_19/A1[12] ),
	.OUT(n2919));
   INVERTER U3312 (.IN(\mult_19/A2[12] ),
	.OUT(n2920));
   INVERTER U3313 (.IN(n2921),
	.OUT(\mult_19/FS_1/PG_int[0][3][0] ));
   INVERTER U3314 (.IN(\mult_19/A2[13] ),
	.OUT(n2922));
   INVERTER U3315 (.IN(n2923),
	.OUT(\mult_19/FS_1/PG_int[0][3][1] ));
   INVERTER U3316 (.IN(\mult_19/FS_1/C[1][3][0] ),
	.OUT(n2924));
   INVERTER U3317 (.IN(\mult_19/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2925));
   INVERTER U3318 (.IN(\mult_19/FS_1/G[1][0][1] ),
	.OUT(n2926));
   INVERTER U3319 (.IN(\mult_19/FS_1/C[1][2][0] ),
	.OUT(n2927));
   INVERTER U3320 (.IN(\mult_19/FS_1/G[1][0][2] ),
	.OUT(n2929));
   INVERTER U3321 (.IN(\mult_19_2/A1[0] ),
	.OUT(n2930));
   INVERTER U3322 (.IN(n2931),
	.OUT(N19));
   INVERTER U3323 (.IN(\mult_19_2/A1[1] ),
	.OUT(n2932));
   INVERTER U3324 (.IN(n2933),
	.OUT(N20));
   INVERTER U3325 (.IN(\mult_19_2/A1[2] ),
	.OUT(n2934));
   INVERTER U3326 (.IN(n2935),
	.OUT(N21));
   INVERTER U3327 (.IN(\mult_19_2/A1[3] ),
	.OUT(n2936));
   INVERTER U3328 (.IN(n2937),
	.OUT(N22));
   INVERTER U3329 (.IN(\mult_19_2/A1[4] ),
	.OUT(n2938));
   INVERTER U3330 (.IN(n2939),
	.OUT(N23));
   INVERTER U3331 (.IN(\mult_19_2/A1[5] ),
	.OUT(n2940));
   INVERTER U3332 (.IN(n2941),
	.OUT(N24));
   INVERTER U3333 (.IN(\mult_19_2/A1[6] ),
	.OUT(n2942));
   INVERTER U3334 (.IN(n2943),
	.OUT(N25));
   INVERTER U3335 (.IN(\mult_19_2/A1[7] ),
	.OUT(n2944));
   INVERTER U3336 (.IN(\mult_19_2/A2[7] ),
	.OUT(n2945));
   INVERTER U3337 (.IN(n2946),
	.OUT(N26));
   INVERTER U3338 (.IN(\mult_19_2/A1[8] ),
	.OUT(n2947));
   INVERTER U3339 (.IN(\mult_19_2/A2[8] ),
	.OUT(n2948));
   INVERTER U3340 (.IN(n2949),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][0] ));
   INVERTER U3341 (.IN(\mult_19_2/A1[9] ),
	.OUT(n2950));
   INVERTER U3342 (.IN(\mult_19_2/A2[9] ),
	.OUT(n2951));
   INVERTER U3343 (.IN(n2952),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][1] ));
   INVERTER U3344 (.IN(n2953),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3345 (.IN(\mult_19_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n2954));
   INVERTER U3346 (.IN(\mult_19_2/A1[10] ),
	.OUT(n2955));
   INVERTER U3347 (.IN(\mult_19_2/A2[10] ),
	.OUT(n2956));
   INVERTER U3348 (.IN(n2957),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][2] ));
   INVERTER U3349 (.IN(n2958),
	.OUT(\mult_19_2/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3350 (.IN(\mult_19_2/FS_1/TEMP_G[0][2][1] ),
	.OUT(n2959));
   INVERTER U3351 (.IN(\mult_19_2/FS_1/C[1][2][1] ),
	.OUT(n2960));
   INVERTER U3352 (.IN(\mult_19_2/FS_1/P[0][2][1] ),
	.OUT(n2961));
   INVERTER U3353 (.IN(\mult_19_2/A1[11] ),
	.OUT(n2962));
   INVERTER U3354 (.IN(\mult_19_2/A2[11] ),
	.OUT(n2963));
   INVERTER U3355 (.IN(n2964),
	.OUT(\mult_19_2/FS_1/PG_int[0][2][3] ));
   INVERTER U3356 (.IN(\mult_19_2/FS_1/TEMP_G[0][2][2] ),
	.OUT(n2965));
   INVERTER U3357 (.IN(\mult_19_2/FS_1/P[0][2][3] ),
	.OUT(n2966));
   INVERTER U3358 (.IN(\mult_19_2/FS_1/C[1][2][2] ),
	.OUT(n2967));
   INVERTER U3359 (.IN(\mult_19_2/FS_1/P[0][2][2] ),
	.OUT(n2968));
   INVERTER U3360 (.IN(\mult_19_2/A1[12] ),
	.OUT(n2969));
   INVERTER U3361 (.IN(\mult_19_2/A2[12] ),
	.OUT(n2970));
   INVERTER U3362 (.IN(n2971),
	.OUT(\mult_19_2/FS_1/PG_int[0][3][0] ));
   INVERTER U3363 (.IN(\mult_19_2/A2[13] ),
	.OUT(n2972));
   INVERTER U3364 (.IN(n2973),
	.OUT(\mult_19_2/FS_1/PG_int[0][3][1] ));
   INVERTER U3365 (.IN(\mult_19_2/FS_1/C[1][3][0] ),
	.OUT(n2974));
   INVERTER U3366 (.IN(\mult_19_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n2975));
   INVERTER U3367 (.IN(\mult_19_2/FS_1/G[1][0][1] ),
	.OUT(n2976));
   INVERTER U3368 (.IN(\mult_19_2/FS_1/C[1][2][0] ),
	.OUT(n2977));
   INVERTER U3369 (.IN(\mult_19_2/FS_1/G[1][0][2] ),
	.OUT(n2979));
   INVERTER U3370 (.IN(\mult_19_3/A1[0] ),
	.OUT(n2980));
   INVERTER U3371 (.IN(n2981),
	.OUT(N51));
   INVERTER U3372 (.IN(\mult_19_3/A1[1] ),
	.OUT(n2982));
   INVERTER U3373 (.IN(n2983),
	.OUT(N52));
   INVERTER U3374 (.IN(\mult_19_3/A1[2] ),
	.OUT(n2984));
   INVERTER U3375 (.IN(n2985),
	.OUT(N53));
   INVERTER U3376 (.IN(\mult_19_3/A1[3] ),
	.OUT(n2986));
   INVERTER U3377 (.IN(n2987),
	.OUT(N54));
   INVERTER U3378 (.IN(\mult_19_3/A1[4] ),
	.OUT(n2988));
   INVERTER U3379 (.IN(n2989),
	.OUT(N55));
   INVERTER U3380 (.IN(\mult_19_3/A1[5] ),
	.OUT(n2990));
   INVERTER U3381 (.IN(n2991),
	.OUT(N56));
   INVERTER U3382 (.IN(\mult_19_3/A1[6] ),
	.OUT(n2992));
   INVERTER U3383 (.IN(n2993),
	.OUT(N57));
   INVERTER U3384 (.IN(\mult_19_3/A1[7] ),
	.OUT(n2994));
   INVERTER U3385 (.IN(\mult_19_3/A2[7] ),
	.OUT(n2995));
   INVERTER U3386 (.IN(n2996),
	.OUT(N58));
   INVERTER U3387 (.IN(\mult_19_3/A1[8] ),
	.OUT(n2997));
   INVERTER U3388 (.IN(\mult_19_3/A2[8] ),
	.OUT(n2998));
   INVERTER U3389 (.IN(n2999),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][0] ));
   INVERTER U3390 (.IN(\mult_19_3/A1[9] ),
	.OUT(n3000));
   INVERTER U3391 (.IN(\mult_19_3/A2[9] ),
	.OUT(n3001));
   INVERTER U3392 (.IN(n3002),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][1] ));
   INVERTER U3393 (.IN(n3003),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3394 (.IN(\mult_19_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3004));
   INVERTER U3395 (.IN(\mult_19_3/A1[10] ),
	.OUT(n3005));
   INVERTER U3396 (.IN(\mult_19_3/A2[10] ),
	.OUT(n3006));
   INVERTER U3397 (.IN(n3007),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][2] ));
   INVERTER U3398 (.IN(n3008),
	.OUT(\mult_19_3/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3399 (.IN(\mult_19_3/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3009));
   INVERTER U3400 (.IN(\mult_19_3/FS_1/C[1][2][1] ),
	.OUT(n3010));
   INVERTER U3401 (.IN(\mult_19_3/FS_1/P[0][2][1] ),
	.OUT(n3011));
   INVERTER U3402 (.IN(\mult_19_3/A1[11] ),
	.OUT(n3012));
   INVERTER U3403 (.IN(\mult_19_3/A2[11] ),
	.OUT(n3013));
   INVERTER U3404 (.IN(n3014),
	.OUT(\mult_19_3/FS_1/PG_int[0][2][3] ));
   INVERTER U3405 (.IN(\mult_19_3/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3015));
   INVERTER U3406 (.IN(\mult_19_3/FS_1/P[0][2][3] ),
	.OUT(n3016));
   INVERTER U3407 (.IN(\mult_19_3/FS_1/C[1][2][2] ),
	.OUT(n3017));
   INVERTER U3408 (.IN(\mult_19_3/FS_1/P[0][2][2] ),
	.OUT(n3018));
   INVERTER U3409 (.IN(\mult_19_3/A1[12] ),
	.OUT(n3019));
   INVERTER U3410 (.IN(\mult_19_3/A2[12] ),
	.OUT(n3020));
   INVERTER U3411 (.IN(n3021),
	.OUT(\mult_19_3/FS_1/PG_int[0][3][0] ));
   INVERTER U3412 (.IN(\mult_19_3/A2[13] ),
	.OUT(n3022));
   INVERTER U3413 (.IN(n3023),
	.OUT(\mult_19_3/FS_1/PG_int[0][3][1] ));
   INVERTER U3414 (.IN(\mult_19_3/FS_1/C[1][3][0] ),
	.OUT(n3024));
   INVERTER U3415 (.IN(\mult_19_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3025));
   INVERTER U3416 (.IN(\mult_19_3/FS_1/G[1][0][1] ),
	.OUT(n3026));
   INVERTER U3417 (.IN(\mult_19_3/FS_1/C[1][2][0] ),
	.OUT(n3027));
   INVERTER U3418 (.IN(\mult_19_3/FS_1/G[1][0][2] ),
	.OUT(n3029));
   INVERTER U3419 (.IN(\mult_20/A1[0] ),
	.OUT(n3030));
   INVERTER U3420 (.IN(n3031),
	.OUT(N83));
   INVERTER U3421 (.IN(\mult_20/A1[1] ),
	.OUT(n3032));
   INVERTER U3422 (.IN(n3033),
	.OUT(N84));
   INVERTER U3423 (.IN(\mult_20/A1[2] ),
	.OUT(n3034));
   INVERTER U3424 (.IN(n3035),
	.OUT(N85));
   INVERTER U3425 (.IN(\mult_20/A1[3] ),
	.OUT(n3036));
   INVERTER U3426 (.IN(n3037),
	.OUT(N86));
   INVERTER U3427 (.IN(\mult_20/A1[4] ),
	.OUT(n3038));
   INVERTER U3428 (.IN(n3039),
	.OUT(N87));
   INVERTER U3429 (.IN(\mult_20/A1[5] ),
	.OUT(n3040));
   INVERTER U3430 (.IN(n3041),
	.OUT(N88));
   INVERTER U3431 (.IN(\mult_20/A1[6] ),
	.OUT(n3042));
   INVERTER U3432 (.IN(n3043),
	.OUT(N89));
   INVERTER U3433 (.IN(\mult_20/A1[7] ),
	.OUT(n3044));
   INVERTER U3434 (.IN(\mult_20/A2[7] ),
	.OUT(n3045));
   INVERTER U3435 (.IN(n3046),
	.OUT(N90));
   INVERTER U3436 (.IN(\mult_20/A1[8] ),
	.OUT(n3047));
   INVERTER U3437 (.IN(\mult_20/A2[8] ),
	.OUT(n3048));
   INVERTER U3438 (.IN(n3049),
	.OUT(\mult_20/FS_1/PG_int[0][2][0] ));
   INVERTER U3439 (.IN(\mult_20/A1[9] ),
	.OUT(n3050));
   INVERTER U3440 (.IN(\mult_20/A2[9] ),
	.OUT(n3051));
   INVERTER U3441 (.IN(n3052),
	.OUT(\mult_20/FS_1/PG_int[0][2][1] ));
   INVERTER U3442 (.IN(n3053),
	.OUT(\mult_20/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3443 (.IN(\mult_20/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3054));
   INVERTER U3444 (.IN(\mult_20/A1[10] ),
	.OUT(n3055));
   INVERTER U3445 (.IN(\mult_20/A2[10] ),
	.OUT(n3056));
   INVERTER U3446 (.IN(n3057),
	.OUT(\mult_20/FS_1/PG_int[0][2][2] ));
   INVERTER U3447 (.IN(n3058),
	.OUT(\mult_20/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3448 (.IN(\mult_20/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3059));
   INVERTER U3449 (.IN(\mult_20/FS_1/C[1][2][1] ),
	.OUT(n3060));
   INVERTER U3450 (.IN(\mult_20/FS_1/P[0][2][1] ),
	.OUT(n3061));
   INVERTER U3451 (.IN(\mult_20/A1[11] ),
	.OUT(n3062));
   INVERTER U3452 (.IN(\mult_20/A2[11] ),
	.OUT(n3063));
   INVERTER U3453 (.IN(n3064),
	.OUT(\mult_20/FS_1/PG_int[0][2][3] ));
   INVERTER U3454 (.IN(\mult_20/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3065));
   INVERTER U3455 (.IN(\mult_20/FS_1/P[0][2][3] ),
	.OUT(n3066));
   INVERTER U3456 (.IN(\mult_20/FS_1/C[1][2][2] ),
	.OUT(n3067));
   INVERTER U3457 (.IN(\mult_20/FS_1/P[0][2][2] ),
	.OUT(n3068));
   INVERTER U3458 (.IN(\mult_20/A1[12] ),
	.OUT(n3069));
   INVERTER U3459 (.IN(\mult_20/A2[12] ),
	.OUT(n3070));
   INVERTER U3460 (.IN(n3071),
	.OUT(\mult_20/FS_1/PG_int[0][3][0] ));
   INVERTER U3461 (.IN(\mult_20/A2[13] ),
	.OUT(n3072));
   INVERTER U3462 (.IN(n3073),
	.OUT(\mult_20/FS_1/PG_int[0][3][1] ));
   INVERTER U3463 (.IN(\mult_20/FS_1/C[1][3][0] ),
	.OUT(n3074));
   INVERTER U3464 (.IN(\mult_20/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3075));
   INVERTER U3465 (.IN(\mult_20/FS_1/G[1][0][1] ),
	.OUT(n3076));
   INVERTER U3466 (.IN(\mult_20/FS_1/C[1][2][0] ),
	.OUT(n3077));
   INVERTER U3467 (.IN(\mult_20/FS_1/G[1][0][2] ),
	.OUT(n3079));
   INVERTER U3468 (.IN(\mult_20_2/A1[0] ),
	.OUT(n3080));
   INVERTER U3469 (.IN(n3081),
	.OUT(N99));
   INVERTER U3470 (.IN(\mult_20_2/A1[1] ),
	.OUT(n3082));
   INVERTER U3471 (.IN(n3083),
	.OUT(N100));
   INVERTER U3472 (.IN(\mult_20_2/A1[2] ),
	.OUT(n3084));
   INVERTER U3473 (.IN(n3085),
	.OUT(N101));
   INVERTER U3474 (.IN(\mult_20_2/A1[3] ),
	.OUT(n3086));
   INVERTER U3475 (.IN(n3087),
	.OUT(N102));
   INVERTER U3476 (.IN(\mult_20_2/A1[4] ),
	.OUT(n3088));
   INVERTER U3477 (.IN(n3089),
	.OUT(N103));
   INVERTER U3478 (.IN(\mult_20_2/A1[5] ),
	.OUT(n3090));
   INVERTER U3479 (.IN(n3091),
	.OUT(N104));
   INVERTER U3480 (.IN(\mult_20_2/A1[6] ),
	.OUT(n3092));
   INVERTER U3481 (.IN(n3093),
	.OUT(N105));
   INVERTER U3482 (.IN(\mult_20_2/A1[7] ),
	.OUT(n3094));
   INVERTER U3483 (.IN(\mult_20_2/A2[7] ),
	.OUT(n3095));
   INVERTER U3484 (.IN(n3096),
	.OUT(N106));
   INVERTER U3485 (.IN(\mult_20_2/A1[8] ),
	.OUT(n3097));
   INVERTER U3486 (.IN(\mult_20_2/A2[8] ),
	.OUT(n3098));
   INVERTER U3487 (.IN(n3099),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][0] ));
   INVERTER U3488 (.IN(\mult_20_2/A1[9] ),
	.OUT(n3100));
   INVERTER U3489 (.IN(\mult_20_2/A2[9] ),
	.OUT(n3101));
   INVERTER U3490 (.IN(n3102),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][1] ));
   INVERTER U3491 (.IN(n3103),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3492 (.IN(\mult_20_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3104));
   INVERTER U3493 (.IN(\mult_20_2/A1[10] ),
	.OUT(n3105));
   INVERTER U3494 (.IN(\mult_20_2/A2[10] ),
	.OUT(n3106));
   INVERTER U3495 (.IN(n3107),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][2] ));
   INVERTER U3496 (.IN(n3108),
	.OUT(\mult_20_2/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3497 (.IN(\mult_20_2/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3109));
   INVERTER U3498 (.IN(\mult_20_2/FS_1/C[1][2][1] ),
	.OUT(n3110));
   INVERTER U3499 (.IN(\mult_20_2/FS_1/P[0][2][1] ),
	.OUT(n3111));
   INVERTER U3500 (.IN(\mult_20_2/A1[11] ),
	.OUT(n3112));
   INVERTER U3501 (.IN(\mult_20_2/A2[11] ),
	.OUT(n3113));
   INVERTER U3502 (.IN(n3114),
	.OUT(\mult_20_2/FS_1/PG_int[0][2][3] ));
   INVERTER U3503 (.IN(\mult_20_2/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3115));
   INVERTER U3504 (.IN(\mult_20_2/FS_1/P[0][2][3] ),
	.OUT(n3116));
   INVERTER U3505 (.IN(\mult_20_2/FS_1/C[1][2][2] ),
	.OUT(n3117));
   INVERTER U3506 (.IN(\mult_20_2/FS_1/P[0][2][2] ),
	.OUT(n3118));
   INVERTER U3507 (.IN(\mult_20_2/A1[12] ),
	.OUT(n3119));
   INVERTER U3508 (.IN(\mult_20_2/A2[12] ),
	.OUT(n3120));
   INVERTER U3509 (.IN(n3121),
	.OUT(\mult_20_2/FS_1/PG_int[0][3][0] ));
   INVERTER U3510 (.IN(\mult_20_2/A2[13] ),
	.OUT(n3122));
   INVERTER U3511 (.IN(n3123),
	.OUT(\mult_20_2/FS_1/PG_int[0][3][1] ));
   INVERTER U3512 (.IN(\mult_20_2/FS_1/C[1][3][0] ),
	.OUT(n3124));
   INVERTER U3513 (.IN(\mult_20_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3125));
   INVERTER U3514 (.IN(\mult_20_2/FS_1/G[1][0][1] ),
	.OUT(n3126));
   INVERTER U3515 (.IN(\mult_20_2/FS_1/C[1][2][0] ),
	.OUT(n3127));
   INVERTER U3516 (.IN(\mult_20_2/FS_1/G[1][0][2] ),
	.OUT(n3129));
   INVERTER U3517 (.IN(\mult_20_3/A1[0] ),
	.OUT(n3130));
   INVERTER U3518 (.IN(n3131),
	.OUT(N131));
   INVERTER U3519 (.IN(\mult_20_3/A1[1] ),
	.OUT(n3132));
   INVERTER U3520 (.IN(n3133),
	.OUT(N132));
   INVERTER U3521 (.IN(\mult_20_3/A1[2] ),
	.OUT(n3134));
   INVERTER U3522 (.IN(n3135),
	.OUT(N133));
   INVERTER U3523 (.IN(\mult_20_3/A1[3] ),
	.OUT(n3136));
   INVERTER U3524 (.IN(n3137),
	.OUT(N134));
   INVERTER U3525 (.IN(\mult_20_3/A1[4] ),
	.OUT(n3138));
   INVERTER U3526 (.IN(n3139),
	.OUT(N135));
   INVERTER U3527 (.IN(\mult_20_3/A1[5] ),
	.OUT(n3140));
   INVERTER U3528 (.IN(n3141),
	.OUT(N136));
   INVERTER U3529 (.IN(\mult_20_3/A1[6] ),
	.OUT(n3142));
   INVERTER U3530 (.IN(n3143),
	.OUT(N137));
   INVERTER U3531 (.IN(\mult_20_3/A1[7] ),
	.OUT(n3144));
   INVERTER U3532 (.IN(\mult_20_3/A2[7] ),
	.OUT(n3145));
   INVERTER U3533 (.IN(n3146),
	.OUT(N138));
   INVERTER U3534 (.IN(\mult_20_3/A1[8] ),
	.OUT(n3147));
   INVERTER U3535 (.IN(\mult_20_3/A2[8] ),
	.OUT(n3148));
   INVERTER U3536 (.IN(n3149),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][0] ));
   INVERTER U3537 (.IN(\mult_20_3/A1[9] ),
	.OUT(n3150));
   INVERTER U3538 (.IN(\mult_20_3/A2[9] ),
	.OUT(n3151));
   INVERTER U3539 (.IN(n3152),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][1] ));
   INVERTER U3540 (.IN(n3153),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3541 (.IN(\mult_20_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3154));
   INVERTER U3542 (.IN(\mult_20_3/A1[10] ),
	.OUT(n3155));
   INVERTER U3543 (.IN(\mult_20_3/A2[10] ),
	.OUT(n3156));
   INVERTER U3544 (.IN(n3157),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][2] ));
   INVERTER U3545 (.IN(n3158),
	.OUT(\mult_20_3/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3546 (.IN(\mult_20_3/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3159));
   INVERTER U3547 (.IN(\mult_20_3/FS_1/C[1][2][1] ),
	.OUT(n3160));
   INVERTER U3548 (.IN(\mult_20_3/FS_1/P[0][2][1] ),
	.OUT(n3161));
   INVERTER U3549 (.IN(\mult_20_3/A1[11] ),
	.OUT(n3162));
   INVERTER U3550 (.IN(\mult_20_3/A2[11] ),
	.OUT(n3163));
   INVERTER U3551 (.IN(n3164),
	.OUT(\mult_20_3/FS_1/PG_int[0][2][3] ));
   INVERTER U3552 (.IN(\mult_20_3/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3165));
   INVERTER U3553 (.IN(\mult_20_3/FS_1/P[0][2][3] ),
	.OUT(n3166));
   INVERTER U3554 (.IN(\mult_20_3/FS_1/C[1][2][2] ),
	.OUT(n3167));
   INVERTER U3555 (.IN(\mult_20_3/FS_1/P[0][2][2] ),
	.OUT(n3168));
   INVERTER U3556 (.IN(\mult_20_3/A1[12] ),
	.OUT(n3169));
   INVERTER U3557 (.IN(\mult_20_3/A2[12] ),
	.OUT(n3170));
   INVERTER U3558 (.IN(n3171),
	.OUT(\mult_20_3/FS_1/PG_int[0][3][0] ));
   INVERTER U3559 (.IN(\mult_20_3/A2[13] ),
	.OUT(n3172));
   INVERTER U3560 (.IN(n3173),
	.OUT(\mult_20_3/FS_1/PG_int[0][3][1] ));
   INVERTER U3561 (.IN(\mult_20_3/FS_1/C[1][3][0] ),
	.OUT(n3174));
   INVERTER U3562 (.IN(\mult_20_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3175));
   INVERTER U3563 (.IN(\mult_20_3/FS_1/G[1][0][1] ),
	.OUT(n3176));
   INVERTER U3564 (.IN(\mult_20_3/FS_1/C[1][2][0] ),
	.OUT(n3177));
   INVERTER U3565 (.IN(\mult_20_3/FS_1/G[1][0][2] ),
	.OUT(n3179));
   INVERTER U3566 (.IN(\mult_21/A1[0] ),
	.OUT(n3180));
   INVERTER U3567 (.IN(n3181),
	.OUT(N163));
   INVERTER U3568 (.IN(\mult_21/A1[1] ),
	.OUT(n3182));
   INVERTER U3569 (.IN(n3183),
	.OUT(N164));
   INVERTER U3570 (.IN(\mult_21/A1[2] ),
	.OUT(n3184));
   INVERTER U3571 (.IN(n3185),
	.OUT(N165));
   INVERTER U3572 (.IN(\mult_21/A1[3] ),
	.OUT(n3186));
   INVERTER U3573 (.IN(n3187),
	.OUT(N166));
   INVERTER U3574 (.IN(\mult_21/A1[4] ),
	.OUT(n3188));
   INVERTER U3575 (.IN(n3189),
	.OUT(N167));
   INVERTER U3576 (.IN(\mult_21/A1[5] ),
	.OUT(n3190));
   INVERTER U3577 (.IN(n3191),
	.OUT(N168));
   INVERTER U3578 (.IN(\mult_21/A1[6] ),
	.OUT(n3192));
   INVERTER U3579 (.IN(n3193),
	.OUT(N169));
   INVERTER U3580 (.IN(\mult_21/A1[7] ),
	.OUT(n3194));
   INVERTER U3581 (.IN(\mult_21/A2[7] ),
	.OUT(n3195));
   INVERTER U3582 (.IN(n3196),
	.OUT(N170));
   INVERTER U3583 (.IN(\mult_21/A1[8] ),
	.OUT(n3197));
   INVERTER U3584 (.IN(\mult_21/A2[8] ),
	.OUT(n3198));
   INVERTER U3585 (.IN(n3199),
	.OUT(\mult_21/FS_1/PG_int[0][2][0] ));
   INVERTER U3586 (.IN(\mult_21/A1[9] ),
	.OUT(n3200));
   INVERTER U3587 (.IN(\mult_21/A2[9] ),
	.OUT(n3201));
   INVERTER U3588 (.IN(n3202),
	.OUT(\mult_21/FS_1/PG_int[0][2][1] ));
   INVERTER U3589 (.IN(n3203),
	.OUT(\mult_21/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3590 (.IN(\mult_21/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3204));
   INVERTER U3591 (.IN(\mult_21/A1[10] ),
	.OUT(n3205));
   INVERTER U3592 (.IN(\mult_21/A2[10] ),
	.OUT(n3206));
   INVERTER U3593 (.IN(n3207),
	.OUT(\mult_21/FS_1/PG_int[0][2][2] ));
   INVERTER U3594 (.IN(n3208),
	.OUT(\mult_21/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3595 (.IN(\mult_21/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3209));
   INVERTER U3596 (.IN(\mult_21/FS_1/C[1][2][1] ),
	.OUT(n3210));
   INVERTER U3597 (.IN(\mult_21/FS_1/P[0][2][1] ),
	.OUT(n3211));
   INVERTER U3598 (.IN(\mult_21/A1[11] ),
	.OUT(n3212));
   INVERTER U3599 (.IN(\mult_21/A2[11] ),
	.OUT(n3213));
   INVERTER U3600 (.IN(n3214),
	.OUT(\mult_21/FS_1/PG_int[0][2][3] ));
   INVERTER U3601 (.IN(\mult_21/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3215));
   INVERTER U3602 (.IN(\mult_21/FS_1/P[0][2][3] ),
	.OUT(n3216));
   INVERTER U3603 (.IN(\mult_21/FS_1/C[1][2][2] ),
	.OUT(n3217));
   INVERTER U3604 (.IN(\mult_21/FS_1/P[0][2][2] ),
	.OUT(n3218));
   INVERTER U3605 (.IN(\mult_21/A1[12] ),
	.OUT(n3219));
   INVERTER U3606 (.IN(\mult_21/A2[12] ),
	.OUT(n3220));
   INVERTER U3607 (.IN(n3221),
	.OUT(\mult_21/FS_1/PG_int[0][3][0] ));
   INVERTER U3608 (.IN(\mult_21/A2[13] ),
	.OUT(n3222));
   INVERTER U3609 (.IN(n3223),
	.OUT(\mult_21/FS_1/PG_int[0][3][1] ));
   INVERTER U3610 (.IN(\mult_21/FS_1/C[1][3][0] ),
	.OUT(n3224));
   INVERTER U3611 (.IN(\mult_21/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3225));
   INVERTER U3612 (.IN(\mult_21/FS_1/G[1][0][1] ),
	.OUT(n3226));
   INVERTER U3613 (.IN(\mult_21/FS_1/C[1][2][0] ),
	.OUT(n3227));
   INVERTER U3614 (.IN(\mult_21/FS_1/G[1][0][2] ),
	.OUT(n3229));
   INVERTER U3615 (.IN(\mult_21_2/A1[0] ),
	.OUT(n3230));
   INVERTER U3616 (.IN(n3231),
	.OUT(N179));
   INVERTER U3617 (.IN(\mult_21_2/A1[1] ),
	.OUT(n3232));
   INVERTER U3618 (.IN(n3233),
	.OUT(N180));
   INVERTER U3619 (.IN(\mult_21_2/A1[2] ),
	.OUT(n3234));
   INVERTER U3620 (.IN(n3235),
	.OUT(N181));
   INVERTER U3621 (.IN(\mult_21_2/A1[3] ),
	.OUT(n3236));
   INVERTER U3622 (.IN(n3237),
	.OUT(N182));
   INVERTER U3623 (.IN(\mult_21_2/A1[4] ),
	.OUT(n3238));
   INVERTER U3624 (.IN(n3239),
	.OUT(N183));
   INVERTER U3625 (.IN(\mult_21_2/A1[5] ),
	.OUT(n3240));
   INVERTER U3626 (.IN(n3241),
	.OUT(N184));
   INVERTER U3627 (.IN(\mult_21_2/A1[6] ),
	.OUT(n3242));
   INVERTER U3628 (.IN(n3243),
	.OUT(N185));
   INVERTER U3629 (.IN(\mult_21_2/A1[7] ),
	.OUT(n3244));
   INVERTER U3630 (.IN(\mult_21_2/A2[7] ),
	.OUT(n3245));
   INVERTER U3631 (.IN(n3246),
	.OUT(N186));
   INVERTER U3632 (.IN(\mult_21_2/A1[8] ),
	.OUT(n3247));
   INVERTER U3633 (.IN(\mult_21_2/A2[8] ),
	.OUT(n3248));
   INVERTER U3634 (.IN(n3249),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][0] ));
   INVERTER U3635 (.IN(\mult_21_2/A1[9] ),
	.OUT(n3250));
   INVERTER U3636 (.IN(\mult_21_2/A2[9] ),
	.OUT(n3251));
   INVERTER U3637 (.IN(n3252),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][1] ));
   INVERTER U3638 (.IN(n3253),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3639 (.IN(\mult_21_2/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3254));
   INVERTER U3640 (.IN(\mult_21_2/A1[10] ),
	.OUT(n3255));
   INVERTER U3641 (.IN(\mult_21_2/A2[10] ),
	.OUT(n3256));
   INVERTER U3642 (.IN(n3257),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][2] ));
   INVERTER U3643 (.IN(n3258),
	.OUT(\mult_21_2/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3644 (.IN(\mult_21_2/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3259));
   INVERTER U3645 (.IN(\mult_21_2/FS_1/C[1][2][1] ),
	.OUT(n3260));
   INVERTER U3646 (.IN(\mult_21_2/FS_1/P[0][2][1] ),
	.OUT(n3261));
   INVERTER U3647 (.IN(\mult_21_2/A1[11] ),
	.OUT(n3262));
   INVERTER U3648 (.IN(\mult_21_2/A2[11] ),
	.OUT(n3263));
   INVERTER U3649 (.IN(n3264),
	.OUT(\mult_21_2/FS_1/PG_int[0][2][3] ));
   INVERTER U3650 (.IN(\mult_21_2/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3265));
   INVERTER U3651 (.IN(\mult_21_2/FS_1/P[0][2][3] ),
	.OUT(n3266));
   INVERTER U3652 (.IN(\mult_21_2/FS_1/C[1][2][2] ),
	.OUT(n3267));
   INVERTER U3653 (.IN(\mult_21_2/FS_1/P[0][2][2] ),
	.OUT(n3268));
   INVERTER U3654 (.IN(\mult_21_2/A1[12] ),
	.OUT(n3269));
   INVERTER U3655 (.IN(\mult_21_2/A2[12] ),
	.OUT(n3270));
   INVERTER U3656 (.IN(n3271),
	.OUT(\mult_21_2/FS_1/PG_int[0][3][0] ));
   INVERTER U3657 (.IN(\mult_21_2/A2[13] ),
	.OUT(n3272));
   INVERTER U3658 (.IN(n3273),
	.OUT(\mult_21_2/FS_1/PG_int[0][3][1] ));
   INVERTER U3659 (.IN(\mult_21_2/FS_1/C[1][3][0] ),
	.OUT(n3274));
   INVERTER U3660 (.IN(\mult_21_2/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3275));
   INVERTER U3661 (.IN(\mult_21_2/FS_1/G[1][0][1] ),
	.OUT(n3276));
   INVERTER U3662 (.IN(\mult_21_2/FS_1/C[1][2][0] ),
	.OUT(n3277));
   INVERTER U3663 (.IN(\mult_21_2/FS_1/G[1][0][2] ),
	.OUT(n3279));
   INVERTER U3664 (.IN(\mult_21_3/A1[0] ),
	.OUT(n3280));
   INVERTER U3665 (.IN(n3281),
	.OUT(N211));
   INVERTER U3666 (.IN(\mult_21_3/A1[1] ),
	.OUT(n3282));
   INVERTER U3667 (.IN(n3283),
	.OUT(N212));
   INVERTER U3668 (.IN(\mult_21_3/A1[2] ),
	.OUT(n3284));
   INVERTER U3669 (.IN(n3285),
	.OUT(N213));
   INVERTER U3670 (.IN(\mult_21_3/A1[3] ),
	.OUT(n3286));
   INVERTER U3671 (.IN(n3287),
	.OUT(N214));
   INVERTER U3672 (.IN(\mult_21_3/A1[4] ),
	.OUT(n3288));
   INVERTER U3673 (.IN(n3289),
	.OUT(N215));
   INVERTER U3674 (.IN(\mult_21_3/A1[5] ),
	.OUT(n3290));
   INVERTER U3675 (.IN(n3291),
	.OUT(N216));
   INVERTER U3676 (.IN(\mult_21_3/A1[6] ),
	.OUT(n3292));
   INVERTER U3677 (.IN(n3293),
	.OUT(N217));
   INVERTER U3678 (.IN(\mult_21_3/A1[7] ),
	.OUT(n3294));
   INVERTER U3679 (.IN(\mult_21_3/A2[7] ),
	.OUT(n3295));
   INVERTER U3680 (.IN(n3296),
	.OUT(N218));
   INVERTER U3681 (.IN(\mult_21_3/A1[8] ),
	.OUT(n3297));
   INVERTER U3682 (.IN(\mult_21_3/A2[8] ),
	.OUT(n3298));
   INVERTER U3683 (.IN(n3299),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][0] ));
   INVERTER U3684 (.IN(\mult_21_3/A1[9] ),
	.OUT(n3300));
   INVERTER U3685 (.IN(\mult_21_3/A2[9] ),
	.OUT(n3301));
   INVERTER U3686 (.IN(n3302),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][1] ));
   INVERTER U3687 (.IN(n3303),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][2][1] ));
   INVERTER U3688 (.IN(\mult_21_3/FS_1/TEMP_P[0][2][0] ),
	.OUT(n3304));
   INVERTER U3689 (.IN(\mult_21_3/A1[10] ),
	.OUT(n3305));
   INVERTER U3690 (.IN(\mult_21_3/A2[10] ),
	.OUT(n3306));
   INVERTER U3691 (.IN(n3307),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][2] ));
   INVERTER U3692 (.IN(n3308),
	.OUT(\mult_21_3/FS_1/TEMP_P[0][2][2] ));
   INVERTER U3693 (.IN(\mult_21_3/FS_1/TEMP_G[0][2][1] ),
	.OUT(n3309));
   INVERTER U3694 (.IN(\mult_21_3/FS_1/C[1][2][1] ),
	.OUT(n3310));
   INVERTER U3695 (.IN(\mult_21_3/FS_1/P[0][2][1] ),
	.OUT(n3311));
   INVERTER U3696 (.IN(\mult_21_3/A1[11] ),
	.OUT(n3312));
   INVERTER U3697 (.IN(\mult_21_3/A2[11] ),
	.OUT(n3313));
   INVERTER U3698 (.IN(n3314),
	.OUT(\mult_21_3/FS_1/PG_int[0][2][3] ));
   INVERTER U3699 (.IN(\mult_21_3/FS_1/TEMP_G[0][2][2] ),
	.OUT(n3315));
   INVERTER U3700 (.IN(\mult_21_3/FS_1/P[0][2][3] ),
	.OUT(n3316));
   INVERTER U3701 (.IN(\mult_21_3/FS_1/C[1][2][2] ),
	.OUT(n3317));
   INVERTER U3702 (.IN(\mult_21_3/FS_1/P[0][2][2] ),
	.OUT(n3318));
   INVERTER U3703 (.IN(\mult_21_3/A1[12] ),
	.OUT(n3319));
   INVERTER U3704 (.IN(\mult_21_3/A2[12] ),
	.OUT(n3320));
   INVERTER U3705 (.IN(n3321),
	.OUT(\mult_21_3/FS_1/PG_int[0][3][0] ));
   INVERTER U3706 (.IN(\mult_21_3/A2[13] ),
	.OUT(n3322));
   INVERTER U3707 (.IN(n3323),
	.OUT(\mult_21_3/FS_1/PG_int[0][3][1] ));
   INVERTER U3708 (.IN(\mult_21_3/FS_1/C[1][3][0] ),
	.OUT(n3324));
   INVERTER U3709 (.IN(\mult_21_3/FS_1/TEMP_P[0][3][0] ),
	.OUT(n3325));
   INVERTER U3710 (.IN(\mult_21_3/FS_1/G[1][0][1] ),
	.OUT(n3326));
   INVERTER U3711 (.IN(\mult_21_3/FS_1/C[1][2][0] ),
	.OUT(n3327));
   INVERTER U3712 (.IN(\mult_21_3/FS_1/G[1][0][2] ),
	.OUT(n3329));
endmodule
