* File: /home/eng/s/sxv240035/cad/gf65/tutorial/MUX21/HSPICE/MUX21.pex.sp
* Created: Tue Dec  3 11:01:01 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "MUX21.pex.sp.pex"
.subckt MUX21  VSS OUT VDD S A B
* 
* B	B
* A	A
* S	S
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=9.75507e-12
+ PERIM=1.2534e-05
XMNMO N_NET11_MNMO_d N_S_MNMO_g N_VSS_MNMO_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.5912e-13 AS=1.17e-13 PD=1.652e-06 PS=9.7e-07
+ NRD=0.196154 NRS=0.413462 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.06e-07 SB=2.313e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.054e-14 PANW9=0 PANW10=0
XMMN1 NET38 N_A_MMN1_g N_VSS_MNMO_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=9.334e-14 AS=1.17e-13 PD=8.79e-07 PS=9.7e-07 NRD=0.345192
+ NRS=0.451923 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07
+ SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.1e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.054e-14 PANW9=0 PANW10=0
XMMN0 N_NET18_MMN0_d N_NET11_MMN0_g NET38 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=8.762e-14 AS=9.334e-14 PD=8.57e-07 PS=8.79e-07 NRD=0.432692
+ NRS=0.345192 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.239e-06
+ SB=1.38e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.1e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.054e-14 PANW9=0 PANW10=0
XMMN2 N_NET18_MMN0_d N_S_MMN2_g NET39 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=8.762e-14 AS=3.666e-14 PD=8.57e-07 PS=6.61e-07 NRD=0.215385
+ NRS=0.135577 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.638e-06
+ SB=9.81e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.1e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.054e-14 PANW9=0 PANW10=0
XMMN3 NET39 N_B_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=3.666e-14 AS=1.0816e-13 PD=6.61e-07 PS=9.36e-07 NRD=0.135577
+ NRS=0.4 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.841e-06 SB=7.78e-07
+ SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.1e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.054e-14 PANW9=0 PANW10=0
XMMN4 N_OUT_MMN4_d N_NET18_MMN4_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.56e-13 AS=1.0816e-13 PD=1.64e-06 PS=9.36e-07
+ NRD=0.309615 NRS=0.4 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=2.319e-06 SB=3e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.054e-14 PANW9=0 PANW10=0
XMMP5 N_NET11_MMP5_d N_S_MMP5_g N_VDD_MMP5_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=2.2032e-13 AS=1.62e-13 PD=2.052e-06 PS=1.17e-06
+ NRD=0.15 NRS=0.440278 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=3.06e-07 SB=2.313e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.728e-15
+ PANW5=3.1e-15 PANW6=4.364e-14 PANW7=1.96e-14 PANW8=1.24e-14 PANW9=7.812e-15
+ PANW10=1.519e-14
XMMP1 NET41 N_A_MMP1_g N_VDD_MMP5_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.2924e-13 AS=1.62e-13 PD=1.079e-06 PS=1.17e-06 NRD=0.249306
+ NRS=0.184722 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07
+ SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.728e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=5.2452e-14 PANW10=1.519e-14
XMMP0 N_NET18_MMP0_d N_S_MMP0_g NET41 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.2132e-13 AS=1.2924e-13 PD=1.057e-06 PS=1.079e-06 NRD=0.313889
+ NRS=0.249306 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.239e-06
+ SB=1.38e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.728e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=7.812e-15 PANW10=1.0447e-13
XMMP2 N_NET18_MMP0_d N_NET11_MMP2_g NET40 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.2132e-13 AS=5.076e-14 PD=1.057e-06 PS=8.61e-07 NRD=0.154167
+ NRS=0.0979167 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.638e-06
+ SB=9.81e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.728e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=7.812e-15 PANW10=1.0447e-13
XMMP3 NET40 N_B_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=5.076e-14 AS=1.4976e-13 PD=8.61e-07 PS=1.136e-06 NRD=0.0979167
+ NRS=0.280556 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.841e-06
+ SB=7.78e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.728e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=5.2452e-14 PANW10=1.519e-14
XMMP4 N_OUT_MMP4_d N_NET18_MMP4_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=2.16e-13 AS=1.4976e-13 PD=2.04e-06 PS=1.136e-06
+ NRD=0.218056 NRS=0.297222 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=2.319e-06 SB=3e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.728e-15
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=3.904e-14 PANW8=3.04e-14 PANW9=7.812e-15
+ PANW10=1.519e-14
*
.include "MUX21.pex.sp.MUX21.pxi"
*
.ends
*
*
