* File: NOR2.pex.sp
* Created: Sun Dec  1 11:28:01 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt NOR2  OUT GND! VDD! A B
* 
XD0_noxref GND! VDD! DIODENWX  AREA=4.95556e-12 PERIM=9.074e-06
XMMN0 OUT A GND! GND! NFET L=6.2e-08 W=7e-07 AD=2.142e-13 AS=1.3615e-13
+ PD=2.012e-06 PS=1.089e-06 NRD=0.194286 NRS=0.275714 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=7.46e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.34e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=1.86e-15
XMMN1 OUT B GND! GND! NFET L=6.2e-08 W=7e-07 AD=2.065e-13 AS=1.3615e-13
+ PD=1.99e-06 PS=1.089e-06 NRD=0.154286 NRS=0.28 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=7.57e-07 SB=2.95e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=4.34e-15 PANW8=1.24e-14 PANW9=2.48e-14 PANW10=1.86e-15
XMMP0 NET16 A VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.5285e-13 AS=3.978e-13
+ PD=1.689e-06 PS=3.212e-06 NRD=0.149615 NRS=0.104615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=7.46e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=7.0576e-14 PANW7=2.54e-14 PANW8=2.1514e-14
+ PANW9=1.302e-13 PANW10=6.5224e-14
XMMP1 OUT B NET16 VDD! PFET L=6.2e-08 W=1.3e-06 AD=3.835e-13 AS=2.5285e-13
+ PD=3.19e-06 PS=1.689e-06 NRD=0.0815385 NRS=0.149615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=7.57e-07 SB=2.95e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=2.976e-15 PANW7=5.01e-14 PANW8=6.5714e-14
+ PANW9=1.289e-13 PANW10=6.5224e-14
*
.include "NOR2.pex.sp.NOR2.pxi"
*
.ends
*
*
