* File: NAND3.pex.sp
* Created: Mon Dec  2 23:31:06 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt NAND3  GND! OUT VDD! C B A
* 
XD0_noxref GND! VDD! DIODENWX  AREA=6.81811e-12 PERIM=1.0484e-05
XMMN0 NET16 C GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.5912e-13
+ PD=9.7e-07 PS=1.652e-06 NRD=0.432692 NRS=0.192308 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMN1 NET17 B NET16 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.432692 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMN2 OUT A NET17 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.5184e-13 AS=1.17e-13
+ PD=1.624e-06 PS=9.7e-07 NRD=0.236538 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMP2 OUT C VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2032e-13
+ PD=1.17e-06 PS=2.052e-06 NRD=0.431944 NRS=0.15 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=3.744e-14 PANW7=7.2e-15 PANW8=9.114e-15 PANW9=3.255e-14
+ PANW10=9.2256e-14
XMMP0 OUT B VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.193056 NRS=0.261111 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=9.114e-15 PANW9=1.2183e-13
+ PANW10=4.7616e-14
XMMP1 OUT A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.1024e-13 AS=1.62e-13
+ PD=2.024e-06 PS=1.17e-06 NRD=0.180556 NRS=0.363889 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=2.88e-14 PANW8=2.4954e-14 PANW9=3.255e-14
+ PANW10=9.2256e-14
*
.include "NAND3.pex.sp.NAND3.pxi"
*
.ends
*
*
