* File: NAND4.pex.sp
* Created: Fri Oct 18 19:15:51 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt NAND4  GND! OUT VDD! D C B A
* 
XD0_noxref GND! VDD! DIODENWX  AREA=8.5004e-12 PERIM=1.169e-05
XMMN3 NET19 D GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=2.142e-13
+ PD=1.15e-06 PS=2.012e-06 NRD=0.321429 NRS=0.142857 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN2 NET20 C NET19 GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.575e-13
+ PD=1.15e-06 PS=1.15e-06 NRD=0.321429 NRS=0.321429 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN1 NET21 B NET20 GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.575e-13
+ PD=1.15e-06 PS=1.15e-06 NRD=0.321429 NRS=0.321429 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN0 OUT A NET21 GND! NFET L=6.2e-08 W=7e-07 AD=2.198e-13 AS=1.575e-13
+ PD=2.028e-06 PS=1.15e-06 NRD=0.175714 NRS=0.321429 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMP3 OUT D VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=3.978e-13
+ PD=1.75e-06 PS=3.212e-06 NRD=0.241538 NRS=0.0830769 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=3.1e-16 PANW6=7.38e-14 PANW7=2.54e-14 PANW8=1.24e-14
+ PANW9=2.9202e-14 PANW10=6.169e-14
XMMP2 OUT C VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=2.925e-13
+ PD=1.75e-06 PS=1.75e-06 NRD=0.104615 NRS=0.241538 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=3.1e-16 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14
+ PANW9=1.09802e-13 PANW10=1.4229e-13
XMMP1 OUT B VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=2.925e-13
+ PD=1.75e-06 PS=1.75e-06 NRD=0.145385 NRS=0.104615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=3.1e-16 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14
+ PANW9=1.09802e-13 PANW10=1.4229e-13
XMMP0 OUT A VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=4.082e-13
+ PD=1.75e-06 PS=3.228e-06 NRD=0.200769 NRS=0.103846 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=3.1e-16 PANW6=3.87e-14 PANW7=6.05e-14 PANW8=1.24e-14
+ PANW9=2.9202e-14 PANW10=6.169e-14
*
.include "NAND4.pex.sp.NAND4.pxi"
*
.ends
*
*
