* File: /home/eng/s/sxv240035/cad/gf65/tutorial/OAI22/HSPICE/OAI22.pex.sp
* Created: Thu Dec  5 19:52:44 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "OAI22.pex.sp.pex"
.subckt OAI22  VSS OUT VDD B D C A
* 
* A	A
* C	C
* D	D
* B	B
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.28285e-11
+ PERIM=1.4672e-05
XMMN0 N_NET12_MMN0_d N_B_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.5912e-13 AS=1.17e-13 PD=1.652e-06 PS=9.7e-07
+ NRD=0.192308 NRS=0.434615 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN1 N_NET12_MMN1_d N_D_MMN1_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.426923
+ NRS=0.430769 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07
+ SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN3 N_OUT_MMN3_d N_C_MMN3_g N_NET12_MMN1_d N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.230769
+ NRS=0.438462 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.33e-06
+ SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN2 N_OUT_MMN3_d N_A_MMN2_g N_NET12_MMN2_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.6328e-13 PD=9.7e-07 PS=1.668e-06 NRD=0.634615
+ NRS=0.223077 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.842e-06
+ SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP3 NET26 N_B_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=2.2032e-13 PD=1.17e-06 PS=2.052e-06 NRD=0.3125
+ NRS=0.15 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=1.85e-06
+ SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
XMMP1 N_OUT_MMP1_d N_D_MMP1_g NET26 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06 NRD=0.330556
+ NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07
+ SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=2.2648e-14
XMMP0 N_OUT_MMP1_d N_C_MMP0_g NET27 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06 NRD=0.294444
+ NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06
+ SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
XMMP2 NET27 N_A_MMP2_g N_VDD_MMP2_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=2.2608e-13 PD=1.17e-06 PS=2.068e-06 NRD=0.3125
+ NRS=0.198611 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.842e-06
+ SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=2.4382e-14 PANW10=4.7848e-14
*
.include "OAI22.pex.sp.OAI22.pxi"
*
.ends
*
*
