* File: Tri_INV.pex.sp
* Created: Fri Oct 18 19:49:12 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt Tri_INV  GND! OUT VDD! EN IN
* 
XD0_noxref GND! VDD! DIODENWX  AREA=7.61944e-12 PERIM=1.1126e-05
XMMN2 NET9 EN GND! GND! NFET L=6.2e-08 W=7e-07 AD=2.142e-13 AS=1.575e-13
+ PD=2.012e-06 PS=1.15e-06 NRD=0.167143 NRS=0.317143 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=2.139e-14 PANW10=2.201e-14
XMMN1 NET15 IN GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.2565e-13 AS=1.575e-13
+ PD=1.059e-06 PS=1.15e-06 NRD=0.274286 NRS=0.325714 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=2.139e-14 PANW10=2.201e-14
XMMN0 OUT EN NET15 GND! NFET L=6.2e-08 W=7e-07 AD=2.681e-13 AS=1.2565e-13
+ PD=2.166e-06 PS=1.059e-06 NRD=0.305714 NRS=0.238571 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.239e-06 SB=3.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=2.139e-14 PANW10=2.201e-14
XMMP2 NET9 EN VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=3.978e-13 AS=2.925e-13
+ PD=3.212e-06 PS=1.75e-06 NRD=0.0830769 NRS=0.241538 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=6.76e-14 PANW7=1.8766e-14 PANW8=1.24e-14
+ PANW9=4.2346e-14 PANW10=1.55e-13
XMMP0 NET15 IN VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.3335e-13 AS=2.925e-13
+ PD=1.659e-06 PS=1.75e-06 NRD=0.145385 NRS=0.104615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=5.766e-15 PANW8=1.24e-14 PANW9=2.03546e-13
+ PANW10=7.44e-14
XMMP1 OUT NET9 NET15 VDD! PFET L=6.2e-08 W=1.3e-06 AD=4.979e-13 AS=2.3335e-13
+ PD=3.366e-06 PS=1.659e-06 NRD=0.173846 NRS=0.130769 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.239e-06 SB=3.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=5.766e-15 PANW8=9.3e-14 PANW9=4.2346e-14
+ PANW10=1.55e-13
*
.include "Tri_INV.pex.sp.TRI_INV.pxi"
*
.ends
*
*
