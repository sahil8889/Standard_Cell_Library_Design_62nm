* File: AOI22.pex.sp
* Created: Mon Dec  2 23:02:32 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt AOI22  GND! OUT VDD! B A C D
* 
XD0_noxref GND! VDD! DIODENWX  AREA=8.18246e-12 PERIM=1.1442e-05
XMMN0 NET25 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.5912e-13
+ PD=9.7e-07 PS=1.652e-06 NRD=0.432692 NRS=0.223077 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14
+ PANW10=0
XMMN2 OUT A NET25 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.405769 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14 PANW10=0
XMMN3 OUT C NET24 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.459615 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14 PANW10=0
XMMN1 NET24 D GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.6328e-13
+ PD=9.7e-07 PS=1.668e-06 NRD=0.432692 NRS=0.225 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=4.774e-15 PANW8=1.24e-14 PANW9=1.5066e-14 PANW10=0
XMMP3 NET26 B VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.2032e-13 AS=1.62e-13
+ PD=2.052e-06 PS=1.17e-06 NRD=0.15 NRS=0.4375 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=3.899e-14 PANW7=1.96e-14 PANW8=1.24e-14 PANW9=1.829e-14
+ PANW10=2.6908e-14
XMMP2 NET26 A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.334722 NRS=0.1875 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=1.55e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=6.293e-14
+ PANW10=7.1548e-14
XMMP0 OUT C NET26 VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.156944 NRS=0.290278 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=1.55e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=6.293e-14
+ PANW10=7.1548e-14
XMMP1 OUT D NET26 VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2608e-13
+ PD=1.17e-06 PS=2.068e-06 NRD=0.468056 NRS=0.197222 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=1.55e-15 PANW7=5.704e-14 PANW8=1.24e-14 PANW9=1.829e-14
+ PANW10=2.6908e-14
c_6 GND! 0 3.8436e-20
c_23 NET26 0 3.8436e-20
*
.include "AOI22.pex.sp.AOI22.pxi"
*
.ends
*
*
