* File: /home/eng/s/sxv240035/cad/gf65/tutorial/XOR2/HSPICE/XOR2.pex.sp
* Created: Thu Dec  5 19:57:34 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "XOR2.pex.sp.pex"
.subckt XOR2  VSS OUT VDD B A
* 
* A	A
* B	B
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.44224e-11
+ PERIM=1.578e-05
XMMN1 N_NET24_MMN1_d N_B_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.0114e-13 AS=1.5912e-13 PD=9.09e-07 PS=1.652e-06
+ NRD=0.361538 NRS=0.261538 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.06e-07 SB=2.271e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN0 N_NET24_MMN1_d N_A_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.0114e-13 AS=1.261e-13 PD=9.09e-07 PS=1.005e-06
+ NRD=0.386538 NRS=0.728846 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=7.57e-07 SB=1.82e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN2 N_OUT_MMN2_d N_NET24_MMN2_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.261e-13 PD=9.7e-07 PS=1.005e-06
+ NRD=0.446154 NRS=0.203846 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.304e-06 SB=1.273e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN4 N_OUT_MMN2_d N_A_MMN4_g NET31 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.17e-13 PD=9.7e-07 PS=9.7e-07 NRD=0.419231
+ NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.816e-06
+ SB=7.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN3 NET31 N_B_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.17e-13 AS=1.2948e-13 PD=9.7e-07 PS=1.538e-06 NRD=0.432692
+ NRS=0.234615 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.328e-06
+ SB=2.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP3 N_NET24_MMP3_d N_B_MMP3_g NET30 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=2.2032e-13 AS=1.4004e-13 PD=2.052e-06 PS=1.109e-06 NRD=0.188889
+ NRS=0.270139 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07
+ SB=2.271e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
XMMP4 NET30 N_A_MMP4_g N_VDD_MMP4_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.4004e-13 AS=1.746e-13 PD=1.109e-06 PS=1.205e-06 NRD=0.270139
+ NRS=0.358333 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.57e-07
+ SB=1.82e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=4.8568e-14
XMMP2 N_NET14_MMP2_d N_NET24_MMP2_g N_VDD_MMP4_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.746e-13 PD=1.17e-06 PS=1.205e-06
+ NRD=0.3125 NRS=0.315278 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.304e-06 SB=1.273e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15
+ PANW10=1.7608e-14
XMMP1 N_OUT_MMP1_d N_A_MMP1_g N_NET14_MMP2_d N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=1.62e-13 PD=1.17e-06 PS=1.17e-06 NRD=0.193056
+ NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.816e-06
+ SB=7.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
XMMP0 N_OUT_MMP1_d N_B_MMP0_g N_NET14_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.62e-13 AS=1.7928e-13 PD=1.17e-06 PS=1.938e-06 NRD=0.431944
+ NRS=0.186111 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.328e-06
+ SB=2.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=6.2248e-14
*
.include "XOR2.pex.sp.XOR2.pxi"
*
.ends
*
*
