* File: XOR2.pex.sp
* Created: Tue Dec  3 02:28:29 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt XOR2  GND! OUT VDD! B A
* 
XD0_noxref GND! VDD! DIODENWX  AREA=9.93119e-12 PERIM=1.263e-05
XMMN1 NET24 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.0114e-13 AS=1.5912e-13
+ PD=9.09e-07 PS=1.652e-06 NRD=0.361538 NRS=0.261538 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=2.271e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.1966e-14 PANW8=1.24e-14 PANW9=7.874e-15
+ PANW10=0
XMMN0 NET24 A GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.0114e-13 AS=1.261e-13
+ PD=9.09e-07 PS=1.005e-06 NRD=0.386538 NRS=0.728846 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=7.57e-07 SB=1.82e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.1966e-14 PANW8=1.24e-14 PANW9=7.874e-15
+ PANW10=0
XMMN2 OUT NET24 GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.261e-13
+ PD=9.7e-07 PS=1.005e-06 NRD=0.446154 NRS=0.203846 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.304e-06 SB=1.273e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.1966e-14 PANW8=1.24e-14 PANW9=7.874e-15
+ PANW10=0
XMMN4 OUT A NET31 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.419231 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=1.816e-06 SB=7.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=1.1966e-14 PANW8=1.24e-14 PANW9=7.874e-15 PANW10=0
XMMN3 NET31 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.2948e-13
+ PD=9.7e-07 PS=1.538e-06 NRD=0.432692 NRS=0.234615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=2.328e-06 SB=2.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.1966e-14 PANW8=1.24e-14 PANW9=7.874e-15
+ PANW10=0
XMMP3 NET24 B NET30 VDD! PFET L=6.2e-08 W=7.2e-07 AD=2.2032e-13 AS=1.4004e-13
+ PD=2.052e-06 PS=1.109e-06 NRD=0.188889 NRS=0.270139 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=2.271e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=3.8184e-14 PANW7=1.96e-14 PANW8=1.24e-14
+ PANW9=1.9096e-14 PANW10=2.1514e-14
XMMP4 NET30 A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.4004e-13 AS=1.746e-13
+ PD=1.109e-06 PS=1.205e-06 NRD=0.270139 NRS=0.358333 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=7.57e-07 SB=1.82e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=7.44e-16 PANW7=1.24e-14 PANW8=1.312e-14 PANW9=6.3016e-14
+ PANW10=2.1514e-14
XMMP2 NET14 NET24 VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.746e-13
+ PD=1.17e-06 PS=1.205e-06 NRD=0.3125 NRS=0.315278 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.304e-06 SB=1.273e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=7.44e-16 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=1.9096e-14
+ PANW10=1.10794e-13
XMMP1 OUT A NET14 VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.193056 NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=1.816e-06 SB=7.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=7.44e-16 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=6.3736e-14
+ PANW10=2.1514e-14
XMMP0 OUT B NET14 VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.7928e-13
+ PD=1.17e-06 PS=1.938e-06 NRD=0.431944 NRS=0.186111 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=2.328e-06 SB=2.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=7.44e-16 PANW7=5.704e-14 PANW8=1.24e-14 PANW9=1.9096e-14
+ PANW10=2.1514e-14
*
.include "XOR2.pex.sp.XOR2.pxi"
*
.ends
*
*
