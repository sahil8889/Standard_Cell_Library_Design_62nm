* File: /home/eng/s/sxv240035/cad/gf65/tutorial/TRI_INV/HSPICE/Tri_INV.pex.sp
* Created: Thu Dec  5 19:54:53 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "Tri_INV.pex.sp.pex"
.subckt TRI_INV  VSS OUT VDD EN IN
* 
* IN	IN
* EN	EN
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.3801e-11
+ PERIM=1.5348e-05
XMMN2 N_NET9_MMN2_d N_EN_MMN2_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.924e-13 AS=1.17e-13 PD=1.78e-06 PS=9.7e-07
+ NRD=0.388462 NRS=0.407692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.7e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN1 N_NET15_MMN1_d N_IN_MMN1_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=9.334e-14 AS=1.17e-13 PD=8.79e-07 PS=9.7e-07
+ NRD=0.365385 NRS=0.457692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=8.82e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN0 N_OUT_MMN0_d N_EN_MMN0_g N_NET15_MMN1_d N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.9916e-13 AS=9.334e-14 PD=1.806e-06 PS=8.79e-07
+ NRD=0.4 NRS=0.325 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.303e-06
+ SB=3.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP2 N_NET9_MMP2_d N_EN_MMP2_g N_VDD_MMP2_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=2.664e-13 AS=1.62e-13 PD=2.18e-06 PS=1.17e-06
+ NRD=0.280556 NRS=0.441667 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=3.7e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15
+ PANW10=6.2248e-14
XMMP0 N_NET15_MMP0_d N_IN_MMP0_g N_VDD_MMP2_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=1.2924e-13 AS=1.62e-13 PD=1.079e-06 PS=1.17e-06
+ NRD=0.261111 NRS=0.183333 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=8.82e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15
+ PANW10=1.7608e-14
XMMP1 N_OUT_MMP1_d N_NET9_MMP1_g N_NET15_MMP0_d N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=2.7576e-13 AS=1.2924e-13 PD=2.206e-06 PS=1.079e-06
+ NRD=0.288889 NRS=0.2375 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.303e-06 SB=3.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15
+ PANW10=3.1288e-14
*
.include "Tri_INV.pex.sp.TRI_INV.pxi"
*
.ends
*
*
