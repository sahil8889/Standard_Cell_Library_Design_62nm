* File: MUX21.pex.sp
* Created: Fri Oct 18 18:51:50 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt MUX21  GND! OUT VDD! S A B
* 
XD0_noxref GND! VDD! DIODENWX  AREA=1.04404e-11 PERIM=1.2932e-05
XMNMO NET11 S GND! GND! NFET L=6.2e-08 W=7e-07 AD=2.142e-13 AS=1.575e-13
+ PD=2.012e-06 PS=1.15e-06 NRD=0.167143 NRS=0.317143 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=2.313e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.24e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=4.96e-15
XMMN1 NET38 A GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.2565e-13 AS=1.575e-13
+ PD=1.059e-06 PS=1.15e-06 NRD=0.256429 NRS=0.325714 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07 SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.24e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=4.96e-15
XMMN0 NET18 NET11 NET38 GND! NFET L=6.2e-08 W=7e-07 AD=1.1795e-13 AS=1.2565e-13
+ PD=1.037e-06 PS=1.059e-06 NRD=0.305714 NRS=0.256429 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.239e-06 SB=1.38e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.24e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=4.96e-15
XMMN2 NET18 S NET39 GND! NFET L=6.2e-08 W=7e-07 AD=1.1795e-13 AS=4.935e-14
+ PD=1.037e-06 PS=8.41e-07 NRD=0.175714 NRS=0.100714 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.638e-06 SB=9.81e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.24e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=4.96e-15
XMMN3 NET39 B GND! GND! NFET L=6.2e-08 W=7e-07 AD=4.935e-14 AS=1.442e-13
+ PD=8.41e-07 PS=1.112e-06 NRD=0.100714 NRS=0.311429 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.841e-06 SB=7.78e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.24e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=4.96e-15
XMMN4 OUT NET18 GND! GND! NFET L=6.2e-08 W=7e-07 AD=2.128e-13 AS=1.442e-13
+ PD=2.008e-06 PS=1.112e-06 NRD=0.251429 NRS=0.277143 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=2.315e-06 SB=3.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.24e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=4.96e-15
XMMP5 NET11 S VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=3.978e-13 AS=2.925e-13
+ PD=3.212e-06 PS=1.75e-06 NRD=0.0830769 NRS=0.241538 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=2.313e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=6.76e-14 PANW7=1.8766e-14 PANW8=1.24e-14
+ PANW9=4.2346e-14 PANW10=7.44e-14
XMMP1 NET41 A VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.3335e-13 AS=2.925e-13
+ PD=1.659e-06 PS=1.75e-06 NRD=0.138077 NRS=0.104615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07 SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=5.766e-15 PANW8=1.24e-14 PANW9=1.22946e-13
+ PANW10=7.44e-14
XMMP0 NET18 S NET41 VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.1905e-13 AS=2.3335e-13
+ PD=1.637e-06 PS=1.659e-06 NRD=0.173846 NRS=0.138077 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.239e-06 SB=1.38e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=5.766e-15 PANW8=1.24e-14 PANW9=4.2346e-14
+ PANW10=2.356e-13
XMMP2 NET18 NET11 NET40 VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.1905e-13 AS=9.165e-14
+ PD=1.637e-06 PS=1.441e-06 NRD=0.0853846 NRS=0.0542308 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.638e-06 SB=9.81e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=5.766e-15 PANW8=1.24e-14 PANW9=4.2346e-14
+ PANW10=2.356e-13
XMMP3 NET40 B VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=9.165e-14 AS=2.678e-13
+ PD=1.441e-06 PS=1.712e-06 NRD=0.0542308 NRS=0.154615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.841e-06 SB=7.78e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=5.766e-15 PANW8=1.24e-14 PANW9=1.22946e-13
+ PANW10=7.44e-14
XMMP4 OUT NET18 VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=3.952e-13 AS=2.678e-13
+ PD=3.208e-06 PS=1.712e-06 NRD=0.130769 NRS=0.162308 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=2.315e-06 SB=3.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=8.6366e-14 PANW8=1.24e-14 PANW9=4.2346e-14
+ PANW10=7.44e-14
*
.include "MUX21.pex.sp.MUX21.pxi"
*
.ends
*
*
