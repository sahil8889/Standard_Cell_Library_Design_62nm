* File: XOR2.pex.sp
* Created: Fri Oct 18 20:02:46 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt XOR2  GND! OUT VDD! B A
* 
XD0_noxref GND! VDD! DIODENWX  AREA=1.02311e-11 PERIM=1.2798e-05
XMMN1 NET24 B GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.3615e-13 AS=1.624e-13
+ PD=1.089e-06 PS=1.864e-06 NRD=0.275714 NRS=0.194286 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=2.32e-07 SB=2.271e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN0 NET24 A GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.3615e-13 AS=1.6975e-13
+ PD=1.089e-06 PS=1.185e-06 NRD=0.28 NRS=0.55 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=6.83e-07 SB=1.82e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN2 OUT NET24 GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.6975e-13
+ PD=1.15e-06 PS=1.185e-06 NRD=0.332857 NRS=0.142857 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.23e-06 SB=1.273e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN4 OUT A NET31 GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.575e-13
+ PD=1.15e-06 PS=1.15e-06 NRD=0.31 NRS=0.321429 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=1.742e-06 SB=7.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN3 NET31 B GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.743e-13
+ PD=1.15e-06 PS=1.898e-06 NRD=0.321429 NRS=0.175714 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=2.254e-06 SB=2.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMP3 NET24 B NET30 VDD! PFET L=6.2e-08 W=1.3e-06 AD=3.016e-13 AS=2.5285e-13
+ PD=3.064e-06 PS=1.689e-06 NRD=0.104615 NRS=0.149615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=2.32e-07 SB=2.271e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=6.76e-14 PANW7=1.3e-14 PANW8=1.0912e-14 PANW9=4.96e-14
+ PANW10=7.44e-14
XMMP4 NET30 A VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.5285e-13 AS=3.1525e-13
+ PD=1.689e-06 PS=1.785e-06 NRD=0.149615 NRS=0.200769 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=6.83e-07 SB=1.82e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=1.2212e-14 PANW9=1.289e-13
+ PANW10=7.44e-14
XMMP2 NET14 NET24 VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=3.1525e-13
+ PD=1.75e-06 PS=1.785e-06 NRD=0.173077 NRS=0.172308 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.23e-06 SB=1.273e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=1.0912e-14 PANW9=4.96e-14
+ PANW10=2.356e-13
XMMP1 OUT A NET14 VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=2.925e-13
+ PD=1.75e-06 PS=1.75e-06 NRD=0.114615 NRS=0.173077 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.742e-06 SB=7.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=1.0912e-14 PANW9=1.302e-13
+ PANW10=7.44e-14
XMMP0 OUT B NET14 VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=3.237e-13
+ PD=1.75e-06 PS=3.098e-06 NRD=0.231538 NRS=0.103846 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=2.254e-06 SB=2.49e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=8.06e-14 PANW8=1.0912e-14 PANW9=4.96e-14
+ PANW10=7.44e-14
*
.include "XOR2.pex.sp.XOR2.pxi"
*
.ends
*
*
