* File: inverter.pex.sp
* Created: Sun Dec  1 11:43:13 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt inverter  GND! OUT VDD! IN
* 
XD0_noxref GND! VDD! DIODENWX  AREA=3.38989e-12 PERIM=7.894e-06
XMMN0 OUT IN GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.862e-13 AS=1.904e-13
+ PD=1.932e-06 PS=1.944e-06 NRD=0.202857 NRS=0.194286 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=2.72e-07 SB=2.66e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.34e-15 PANW8=1.24e-14 PANW9=2.48e-14
+ PANW10=1.86e-15
XMMP0 OUT IN VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=3.458e-13 AS=3.536e-13
+ PD=3.132e-06 PS=3.144e-06 NRD=0.101538 NRS=0.104615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=2.72e-07 SB=2.66e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=7.1878e-14 PANW7=1.06e-13 PANW8=2.1514e-14
+ PANW9=4.96e-14 PANW10=6.3922e-14
*
.include "inverter.pex.sp.INVERTER.pxi"
*
.ends
*
*
