* File: /home/eng/s/sxv240035/cad/gf65/lib_cell/NOR3/NOR3_LVS/NOR3.pex.sp
* Created: Sat Oct 19 23:51:38 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt NOR3  GND! OUT VDD! A B C
* 
XD0_noxref GND! VDD! DIODENWX  AREA=6.96652e-12 PERIM=1.0708e-05
XMMN1 OUT A GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=2.142e-13
+ PD=1.15e-06 PS=2.012e-06 NRD=0.455714 NRS=0.142857 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN0 OUT B GND! GND! NFET L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.575e-13
+ PD=1.15e-06 PS=1.15e-06 NRD=0.187143 NRS=0.264286 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN2 OUT C GND! GND! NFET L=6.2e-08 W=7e-07 AD=2.044e-13 AS=1.575e-13
+ PD=1.984e-06 PS=1.15e-06 NRD=0.175714 NRS=0.378571 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMP2 NET20 A VDD! VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=3.978e-13
+ PD=1.75e-06 PS=3.212e-06 NRD=0.173077 NRS=0.0830769 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=3.1e-16 PANW6=7.38e-14 PANW7=2.54e-14 PANW8=1.24e-14
+ PANW9=2.9202e-14 PANW10=1.4229e-13
XMMP1 NET21 B NET20 VDD! PFET L=6.2e-08 W=1.3e-06 AD=2.925e-13 AS=2.925e-13
+ PD=1.75e-06 PS=1.75e-06 NRD=0.173077 NRS=0.173077 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=3.1e-16 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14
+ PANW9=1.90402e-13 PANW10=6.169e-14
XMMP0 OUT C NET21 VDD! PFET L=6.2e-08 W=1.3e-06 AD=3.796e-13 AS=2.925e-13
+ PD=3.184e-06 PS=1.75e-06 NRD=0.103846 NRS=0.173077 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=3.1e-16 PANW6=1.14e-14 PANW7=8.78e-14 PANW8=1.24e-14
+ PANW9=2.9202e-14 PANW10=1.4229e-13
*
.include "/home/eng/s/sxv240035/cad/gf65/lib_cell/NOR3/NOR3_LVS/NOR3.pex.sp.NOR3.pxi"
*
.ends
*
*
