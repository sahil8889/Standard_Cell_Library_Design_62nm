* File: /home/eng/s/sxv240035/cad/gf65/tutorial/NOR2/HSPICE/NOR2.pex.sp
* Created: Thu Dec  5 19:46:34 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "NOR2.pex.sp.pex"
.subckt NOR2  OUT VSS VDD A B
* 
* B	B
* A	A
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.00148e-11
+ PERIM=1.2716e-05
XMMN0 N_OUT_MMN0_d N_A_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.5912e-13 AS=1.0114e-13 PD=1.652e-06 PS=9.09e-07 NRD=0.261538
+ NRS=0.359615 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07
+ SB=7.46e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN1 N_OUT_MMN1_d N_B_MMN1_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.534e-13 AS=1.0114e-13 PD=1.63e-06 PS=9.09e-07 NRD=0.215385
+ NRS=0.388462 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=7.57e-07
+ SB=2.95e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP0 NET16 N_A_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.4004e-13 AS=2.2032e-13 PD=1.109e-06 PS=2.052e-06 NRD=0.270139
+ NRS=0.188889 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07
+ SB=7.46e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.06888e-13
XMMP1 N_OUT_MMP1_d N_B_MMP1_g NET16 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=2.124e-13 AS=1.4004e-13 PD=2.03e-06 PS=1.109e-06 NRD=0.155556
+ NRS=0.270139 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.57e-07
+ SB=2.95e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=3.8782e-14 PANW10=3.3448e-14
*
.include "NOR2.pex.sp.NOR2.pxi"
*
.ends
*
*
