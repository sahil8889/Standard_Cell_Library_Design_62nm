* File: OAI21.pex.sp
* Created: Tue Dec  3 01:05:41 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt OAI21  GND! OUT VDD! A B C
* 
XD0_noxref GND! VDD! DIODENWX  AREA=6.79365e-12 PERIM=1.0494e-05
XMMN NET014 A GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.5912e-13 AS=1.17e-13
+ PD=1.652e-06 PS=9.7e-07 NRD=0.192308 NRS=0.605769 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMN0 NET014 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.361538 NRS=0.259615 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMN1 OUT C NET014 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.5184e-13 AS=1.17e-13
+ PD=1.624e-06 PS=9.7e-07 NRD=0.259615 NRS=0.503846 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMP1 NET19 A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2032e-13
+ PD=1.17e-06 PS=2.052e-06 NRD=0.3125 NRS=0.15 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=3.06e-07 SB=1.316e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=3.744e-14 PANW7=7.2e-15 PANW8=9.114e-15 PANW9=2.7962e-14
+ PANW10=9.2566e-14
XMMP0 OUT B NET19 VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.302778 NRS=0.3125 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=8.18e-07 SB=8.04e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=9.114e-15 PANW9=1.17242e-13 PANW10=4.7926e-14
XMMP2 OUT C VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.1024e-13
+ PD=1.17e-06 PS=2.024e-06 NRD=0.322222 NRS=0.191667 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06 SB=2.92e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.464e-14 PANW8=9.114e-15 PANW9=2.7962e-14
+ PANW10=9.2566e-14
c_6 NET014 0 2.79161e-20
c_22 VDD! 0 2.79161e-20
*
.include "OAI21.pex.sp.OAI21.pxi"
*
.ends
*
*
