* File: MUX21.pex.sp
* Created: Sun Dec  1 23:51:02 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt MUX21  GND! OUT VDD! S A B
* 
XD0_noxref GND! VDD! DIODENWX  AREA=8.55304e-12 PERIM=1.1824e-05
XMNMO NET11 S GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.5912e-13 AS=1.17e-13
+ PD=1.652e-06 PS=9.7e-07 NRD=0.225 NRS=0.405769 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=3.06e-07 SB=2.313e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=1.0044e-14 PANW8=1.24e-14 PANW9=9.796e-15 PANW10=0
XMMN1 NET38 A GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=9.334e-14 AS=1.17e-13
+ PD=8.79e-07 PS=9.7e-07 NRD=0.345192 NRS=0.459615 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=8.18e-07 SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.0044e-14 PANW8=1.24e-14 PANW9=9.796e-15
+ PANW10=0
XMMN0 NET18 NET11 NET38 GND! NFET L=6.2e-08 W=5.2e-07 AD=8.762e-14 AS=9.334e-14
+ PD=8.57e-07 PS=8.79e-07 NRD=0.442308 NRS=0.345192 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.239e-06 SB=1.38e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.0044e-14 PANW8=1.24e-14 PANW9=9.796e-15
+ PANW10=0
XMMN2 NET18 S NET39 GND! NFET L=6.2e-08 W=5.2e-07 AD=8.762e-14 AS=3.666e-14
+ PD=8.57e-07 PS=6.61e-07 NRD=0.205769 NRS=0.135577 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.638e-06 SB=9.81e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.0044e-14 PANW8=1.24e-14 PANW9=9.796e-15
+ PANW10=0
XMMN3 NET39 B GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=3.666e-14 AS=1.0816e-13
+ PD=6.61e-07 PS=9.36e-07 NRD=0.135577 NRS=0.403846 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.841e-06 SB=7.78e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.0044e-14 PANW8=1.24e-14 PANW9=9.796e-15
+ PANW10=0
XMMN4 OUT NET18 GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.56e-13 AS=1.0816e-13
+ PD=1.64e-06 PS=9.36e-07 NRD=0.311538 NRS=0.396154 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=2.319e-06 SB=3e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=1.0044e-14 PANW8=1.24e-14 PANW9=9.796e-15
+ PANW10=0
XMMP5 NET11 S VDD! VDD! PFET L=6.2e-08 W=7.96e-07 AD=2.43576e-13 AS=1.791e-13
+ PD=2.204e-06 PS=1.246e-06 NRD=0.135678 NRS=0.395729 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07 SB=2.313e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=2.728e-15 PANW5=3.1e-15 PANW6=4.7592e-14 PANW7=2.036e-14 PANW8=1.24e-14
+ PANW9=1.7236e-14 PANW10=3.72e-14
XMMP1 NET41 A VDD! VDD! PFET L=6.2e-08 W=7.96e-07 AD=1.42882e-13 AS=1.791e-13
+ PD=1.155e-06 PS=1.246e-06 NRD=0.225503 NRS=0.169598 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07 SB=1.801e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=2.728e-15 PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14
+ PANW9=6.6588e-14 PANW10=3.72e-14
XMMP0 NET18 S NET41 VDD! PFET L=6.2e-08 W=7.96e-07 AD=1.34126e-13 AS=1.42882e-13
+ PD=1.133e-06 PS=1.155e-06 NRD=0.287688 NRS=0.225503 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.239e-06 SB=1.38e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=2.728e-15 PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14
+ PANW9=1.7236e-14 PANW10=1.35904e-13
XMMP2 NET18 NET11 NET40 VDD! PFET L=6.2e-08 W=7.96e-07 AD=1.34126e-13
+ AS=5.6118e-14 PD=1.133e-06 PS=9.37e-07 NRD=0.135678 NRS=0.0885678 M=1 NF=1
+ CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.638e-06 SB=9.81e-07 SD=0 PANW1=0
+ PANW2=0 PANW3=0 PANW4=2.728e-15 PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14
+ PANW8=1.24e-14 PANW9=1.7236e-14 PANW10=1.35904e-13
XMMP3 NET40 B VDD! VDD! PFET L=6.2e-08 W=7.96e-07 AD=5.6118e-14 AS=1.65568e-13
+ PD=9.37e-07 PS=1.212e-06 NRD=0.0885678 NRS=0.252513 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.841e-06 SB=7.78e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=2.728e-15 PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14
+ PANW9=6.6588e-14 PANW10=3.72e-14
XMMP4 OUT NET18 VDD! VDD! PFET L=6.2e-08 W=7.96e-07 AD=2.388e-13 AS=1.65568e-13
+ PD=2.192e-06 PS=1.212e-06 NRD=0.208543 NRS=0.270101 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=2.319e-06 SB=3e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=2.728e-15 PANW5=3.1e-15 PANW6=6.2e-15 PANW7=4.1852e-14 PANW8=3.23e-14
+ PANW9=1.7236e-14 PANW10=3.72e-14
*
.include "MUX21.pex.sp.MUX21.pxi"
*
.ends
*
*
