* File: /home/eng/s/sxv240035/cad/gf65/lib_cell/OAI22/HSPICE/OAI22.pex.sp
* Created: Thu Oct 24 16:10:19 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "/home/eng/s/sxv240035/cad/gf65/lib_cell/OAI22/HSPICE/OAI22.pex.sp.pex"
.subckt OAI22  GND! OUT VDD! B D C A
* 
* A	A
* C	C
* D	D
* B	B
* VDD!	VDD!
* OUT	OUT
* GND!	GND!
XD0_noxref N_GND!_D0_noxref_pos N_VDD!_D0_noxref_neg DIODENWX  AREA=8.5004e-12
+ PERIM=1.169e-05
XMMN0 N_NET12_MMN0_d N_B_MMN0_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET
+ L=6.2e-08 W=7e-07 AD=2.142e-13 AS=1.575e-13 PD=2.012e-06 PS=1.15e-06
+ NRD=0.142857 NRS=0.328571 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN1 N_NET12_MMN1_d N_D_MMN1_g N_GND!_MMN0_s N_GND!_D0_noxref_pos NFET
+ L=6.2e-08 W=7e-07 AD=1.575e-13 AS=1.575e-13 PD=1.15e-06 PS=1.15e-06
+ NRD=0.315714 NRS=0.314286 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=0 PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN3 N_OUT_MMN3_d N_C_MMN3_g N_NET12_MMN1_d N_GND!_D0_noxref_pos NFET L=6.2e-08
+ W=7e-07 AD=1.575e-13 AS=1.575e-13 PD=1.15e-06 PS=1.15e-06 NRD=0.142857
+ NRS=0.327143 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.33e-06
+ SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMN2 N_OUT_MMN3_d N_A_MMN2_g N_NET12_MMN2_s N_GND!_D0_noxref_pos NFET L=6.2e-08
+ W=7e-07 AD=1.575e-13 AS=2.198e-13 PD=1.15e-06 PS=2.028e-06 NRD=0.5
+ NRS=0.175714 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.842e-06
+ SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=0 PANW9=1.2028e-14 PANW10=3.1372e-14
XMMP3 NET26 N_B_MMP3_g N_VDD!_MMP3_s N_VDD!_D0_noxref_neg PFET L=6.2e-08
+ W=1.3e-06 AD=2.925e-13 AS=3.978e-13 PD=1.75e-06 PS=3.212e-06 NRD=0.173077
+ NRS=0.0830769 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07
+ SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=6.76e-14
+ PANW7=1.3e-14 PANW8=1.0912e-14 PANW9=4.96e-14 PANW10=7.44e-14
XMMP1 N_OUT_MMP1_d N_D_MMP1_g NET26 N_VDD!_D0_noxref_neg PFET L=6.2e-08
+ W=1.3e-06 AD=2.925e-13 AS=2.925e-13 PD=1.75e-06 PS=1.75e-06 NRD=0.182308
+ NRS=0.173077 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=8.18e-07
+ SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=1.0912e-14 PANW9=1.302e-13 PANW10=1.55e-13
XMMP0 N_OUT_MMP1_d N_C_MMP0_g NET27 N_VDD!_D0_noxref_neg PFET L=6.2e-08
+ W=1.3e-06 AD=2.925e-13 AS=2.925e-13 PD=1.75e-06 PS=1.75e-06 NRD=0.163846
+ NRS=0.173077 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06
+ SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=0
+ PANW8=1.0912e-14 PANW9=1.302e-13 PANW10=1.55e-13
XMMP2 NET27 N_A_MMP2_g N_VDD!_MMP2_s N_VDD!_D0_noxref_neg PFET L=6.2e-08
+ W=1.3e-06 AD=2.925e-13 AS=4.082e-13 PD=1.75e-06 PS=3.228e-06 NRD=0.173077
+ NRS=0.103846 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.842e-06
+ SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=3.25e-14
+ PANW7=4.81e-14 PANW8=1.0912e-14 PANW9=4.96e-14 PANW10=7.44e-14
*
.include "/home/eng/s/sxv240035/cad/gf65/lib_cell/OAI22/HSPICE/OAI22.pex.sp.OAI22.pxi"
*
.ends
*
*
