* File: /home/eng/s/sxv240035/cad/gf65/tutorial/NAND2/HSPICE/NAND2.pex.sp
* Created: Thu Dec  5 19:35:18 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "NAND2.pex.sp.pex"
.subckt NAND2  VSS OUT VDD B A
* 
* A	A
* B	B
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.0783e-11
+ PERIM=1.325e-05
XMMN1 NET16 N_B_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.0114e-13 AS=1.5912e-13 PD=9.09e-07 PS=1.652e-06 NRD=0.374038
+ NRS=0.261538 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07
+ SB=7.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN0 N_OUT_MMN0_d N_A_MMN0_g NET16 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=1.43e-13 AS=1.0114e-13 PD=1.59e-06 PS=9.09e-07 NRD=0.217308
+ NRS=0.374038 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=7.57e-07
+ SB=2.75e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP0 N_OUT_MMP0_d N_B_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=2.2032e-13 AS=1.4004e-13 PD=2.052e-06 PS=1.109e-06 NRD=0.188889
+ NRS=0.258333 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.06e-07
+ SB=7.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.418e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.122e-15 PANW10=1.04308e-13
XMMP1 N_OUT_MMP1_d N_A_MMP1_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.98e-13 AS=1.4004e-13 PD=1.99e-06 PS=1.109e-06 NRD=0.156944
+ NRS=0.281944 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.57e-07
+ SB=2.75e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.418e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.122e-15 PANW10=6.0388e-14
*
.include "NAND2.pex.sp.NAND2.pxi"
*
.ends
*
*
