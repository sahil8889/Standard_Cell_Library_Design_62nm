* File: /home/eng/s/sxv240035/cad/gf65/tutorial/DFF/hspice/dff.pex.sp
* Created: Thu Dec  5 19:29:28 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "dff.pex.sp.pex"
.subckt DFF  VSS CLK Q VDD D R
* 
* R	R
* D	D
* VDD	VDD
* Q	Q
* CLK	CLK
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=2.57866e-11
+ PERIM=2.368e-05
XMMN4 NET56 N_D_MMN4_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=3.38e-14 AS=8.32e-14 PD=6.5e-07 PS=1.36e-06 NRD=0.125
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.6e-07
+ SB=1.429e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN3 N_A_MMN3_d N_CLK_MMN3_g NET56 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=5.2e-14 AS=3.38e-14 PD=7.2e-07 PS=6.5e-07 NRD=0.192308 NRS=0.125
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.52e-07 SB=1.237e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=1.1036e-14
+ PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN7 N_A_MMN3_d N_!CLK_MMN7_g NET058 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=5.2e-14 AS=3.38e-14 PD=7.2e-07 PS=6.5e-07 NRD=0.192308 NRS=0.125
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=6.14e-07 SB=9.75e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=1.1036e-14
+ PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN8 NET058 N_B_MMN8_g N_VSS_MMN8_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=3.38e-14 AS=7.748e-14 PD=6.5e-07 PS=8.18e-07 NRD=0.125
+ NRS=0.380769 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=8.06e-07
+ SB=7.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP6 N_B_MMP6_d N_R_MMP6_g N_VSS_MMN8_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=5.226e-14 AS=7.748e-14 PD=7.21e-07 PS=8.18e-07 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.166e-06
+ SB=4.23e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP5 N_B_MMP6_d N_A_MMP5_g N_VSS_MMP5_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=5.226e-14 AS=8.32e-14 PD=7.21e-07 PS=1.36e-06 NRD=0.194231
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.429e-06
+ SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN2 N_!CLK_MMN2_d N_CLK_MMN2_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=8.372e-14 AS=1.1388e-13 PD=1.362e-06 PS=9.58e-07
+ NRD=0.192308 NRS=0.65 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.61e-07 SB=7.77e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN1 N_CLK_MMN1_d N_!CLK_MMN1_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.4404e-13 AS=1.1388e-13 PD=1.594e-06 PS=9.58e-07
+ NRD=0.192308 NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=6.61e-07 SB=2.77e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN15 N_Q_MMN15_d N_C_MMN15_g N_VSS_MMN15_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=1.352e-13 AS=6.76e-14 PD=1.56e-06 PS=7.8e-07
+ NRD=0.384615 NRS=0.307692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=2.6e-07 SB=1.774e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN10 NET057 N_B_MMN10_g N_VSS_MMN15_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=3.38e-14 AS=6.76e-14 PD=6.5e-07 PS=7.8e-07 NRD=0.125 NRS=0.192308
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=5.82e-07 SB=1.452e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=1.1036e-14
+ PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN9 N_C_MMN9_d N_!CLK_MMN9_g NET057 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=5.2e-14 AS=3.38e-14 PD=7.2e-07 PS=6.5e-07 NRD=0.192308 NRS=0.125
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=7.74e-07 SB=1.26e-06 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=1.1036e-14
+ PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN13 N_C_MMN9_d N_CLK_MMN13_g NET056 N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=5.2e-14 AS=3.38e-14 PD=7.2e-07 PS=6.5e-07 NRD=0.192308 NRS=0.125
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.036e-06 SB=9.98e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=1.1036e-14
+ PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN14 NET056 N_E_MMN14_g N_VSS_MMN14_s N_VSS_D0_noxref_pos NFET L=6.2e-08
+ W=5.2e-07 AD=3.38e-14 AS=6.76e-14 PD=6.5e-07 PS=7.8e-07 NRD=0.125 NRS=0.307692
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.228e-06 SB=8.06e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0 PANW7=1.1036e-14
+ PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN12 N_E_MMN12_d N_R_MMN12_g N_VSS_MMN14_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=6.812e-14 AS=6.76e-14 PD=7.82e-07 PS=7.8e-07
+ NRD=0.311538 NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.55e-06 SB=4.84e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMN11 N_E_MMN12_d N_C_MMN11_g N_VSS_MMN11_s N_VSS_D0_noxref_pos NFET
+ L=6.2e-08 W=5.2e-07 AD=6.812e-14 AS=8.32e-14 PD=7.82e-07 PS=1.36e-06
+ NRD=0.192308 NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.874e-06 SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0 PANW5=0 PANW6=0
+ PANW7=1.1036e-14 PANW8=1.24e-14 PANW9=8.804e-15 PANW10=0
XMMP4 NET51 N_D_MMP4_g N_VDD_MMP4_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=4.68e-14 AS=1.152e-13 PD=8.5e-07 PS=1.76e-06 NRD=0.0902778
+ NRS=0.138889 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.6e-07
+ SB=1.429e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.7608e-14
XMMP3 N_A_MMP3_d N_!CLK_MMP3_g NET51 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=7.2e-14 AS=4.68e-14 PD=9.2e-07 PS=8.5e-07 NRD=0.138889
+ NRS=0.0902778 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.52e-07
+ SB=1.237e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.7608e-14
XMMP7 N_A_MMP3_d N_CLK_MMP7_g NET053 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=7.2e-14 AS=4.68e-14 PD=9.2e-07 PS=8.5e-07 NRD=0.138889
+ NRS=0.0902778 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=6.14e-07
+ SB=9.75e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.7608e-14
XMMP8 NET053 N_B_MMP8_g N_VDD_MMP8_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=4.68e-14 AS=1.0728e-13 PD=8.5e-07 PS=1.018e-06 NRD=0.0902778
+ NRS=0.215278 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1 SA=8.06e-07
+ SB=7.83e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.7608e-14
XMMN6 NET58 N_R_MMN6_g N_VDD_MMP8_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=7.236e-14 AS=1.0728e-13 PD=9.21e-07 PS=1.018e-06 NRD=0.139583
+ NRS=0.198611 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.166e-06
+ SB=4.23e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.7608e-14
XMMN5 N_B_MMN5_d N_A_MMN5_g NET58 N_VDD_D0_noxref_neg PFET L=6.2e-08 W=7.2e-07
+ AD=1.152e-13 AS=7.236e-14 PD=1.76e-06 PS=9.21e-07 NRD=0.138889 NRS=0.139583
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.429e-06 SB=1.6e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=0 PANW4=5.58e-16 PANW5=3.1e-15 PANW6=6.2e-15
+ PANW7=1.24e-14 PANW8=1.24e-14 PANW9=9.982e-15 PANW10=1.7608e-14
XMMP2 N_!CLK_MMP2_d N_CLK_MMP2_g N_VDD_MMP2_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=1.1592e-13 AS=1.5768e-13 PD=1.762e-06 PS=1.158e-06
+ NRD=0.138889 NRS=0.254167 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.61e-07 SB=7.77e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15
+ PANW10=1.5686e-14
XMMP1 N_CLK_MMP1_d N_!CLK_MMP1_g N_VDD_MMP2_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=1.9944e-13 AS=1.5768e-13 PD=1.994e-06 PS=1.158e-06
+ NRD=0.138889 NRS=0.354167 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=6.61e-07 SB=2.77e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15
+ PANW10=1.5686e-14
XMMP15 N_Q_MMP15_d N_C_MMP15_g N_VDD_MMP15_s N_VDD_D0_noxref_neg PFET
+ L=6.2e-08 W=7.2e-07 AD=1.872e-13 AS=9.36e-14 PD=1.96e-06 PS=9.8e-07
+ NRD=0.277778 NRS=0.222222 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1
+ SA=2.6e-07 SB=1.774e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15
+ PANW5=3.1e-15 PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15
+ PANW10=1.5686e-14
XMMP10 NET052 N_B_MMP10_g N_VDD_MMP15_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=4.68e-14 AS=9.36e-14 PD=8.5e-07 PS=9.8e-07 NRD=0.0902778
+ NRS=0.138889 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=5.82e-07
+ SB=1.452e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15 PANW10=1.5686e-14
XMMP9 N_C_MMP9_d N_CLK_MMP9_g NET052 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=7.2e-14 AS=4.68e-14 PD=9.2e-07 PS=8.5e-07 NRD=0.138889
+ NRS=0.0902778 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.74e-07
+ SB=1.26e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15 PANW10=1.5686e-14
XMMP13 N_C_MMP9_d N_!CLK_MMP13_g NET050 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=7.2e-14 AS=4.68e-14 PD=9.2e-07 PS=8.5e-07 NRD=0.138889
+ NRS=0.0902778 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.036e-06
+ SB=9.98e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15 PANW10=1.5686e-14
XMMP14 NET050 N_E_MMP14_g N_VDD_MMP14_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=4.68e-14 AS=9.36e-14 PD=8.5e-07 PS=9.8e-07 NRD=0.0902778
+ NRS=0.222222 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1 SA=1.228e-06
+ SB=8.06e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15 PANW10=1.5686e-14
XMMP12 NET051 N_R_MMP12_g N_VDD_MMP14_s N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=9.432e-14 AS=9.36e-14 PD=9.82e-07 PS=9.8e-07 NRD=0.181944
+ NRS=0.138889 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.55e-06
+ SB=4.84e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15 PANW10=1.5686e-14
XMMP11 N_E_MMP11_d N_C_MMP11_g NET051 N_VDD_D0_noxref_neg PFET L=6.2e-08
+ W=7.2e-07 AD=1.152e-13 AS=9.432e-14 PD=1.76e-06 PS=9.82e-07 NRD=0.138889
+ NRS=0.181944 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.874e-06
+ SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=2.48e-15 PANW5=3.1e-15
+ PANW6=6.2e-15 PANW7=1.24e-14 PANW8=1.24e-14 PANW9=8.06e-15 PANW10=6.0326e-14
*
.include "dff.pex.sp.DFF.pxi"
*
.ends
*
*
