* File: NAND4.pex.sp
* Created: Tue Dec  3 00:06:08 2024
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.subckt NAND4  GND! OUT VDD! D C B A
* 
XD0_noxref GND! VDD! DIODENWX  AREA=8.05705e-12 PERIM=1.1354e-05
XMMN3 NET19 D GND! GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.5912e-13
+ PD=9.7e-07 PS=1.652e-06 NRD=0.432692 NRS=0.192308 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMN2 NET20 C NET19 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.432692 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMN1 NET21 B NET20 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.17e-13 AS=1.17e-13
+ PD=9.7e-07 PS=9.7e-07 NRD=0.432692 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=0 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMN0 OUT A NET21 GND! NFET L=6.2e-08 W=5.2e-07 AD=1.6328e-13 AS=1.17e-13
+ PD=1.668e-06 PS=9.7e-07 NRD=0.255769 NRS=0.432692 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=0 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=5.58e-15 PANW9=2.48e-14 PANW10=1.86e-15
XMMP3 OUT D VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2032e-13
+ PD=1.17e-06 PS=2.052e-06 NRD=0.4375 NRS=0.15 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=3.06e-07 SB=1.85e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=3.744e-14 PANW7=7.2e-15 PANW8=9.114e-15 PANW9=3.348e-14
+ PANW10=4.6686e-14
XMMP2 OUT C VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.1875 NRS=0.436111 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0
+ PAR=1 PTWELL=1 SA=8.18e-07 SB=1.338e-06 SD=0 PANW1=0 PANW2=0 PANW3=0 PANW4=0
+ PANW5=0 PANW6=0 PANW7=0 PANW8=9.114e-15 PANW9=7.812e-14 PANW10=9.1326e-14
XMMP1 OUT B VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=1.62e-13
+ PD=1.17e-06 PS=1.17e-06 NRD=0.255556 NRS=0.188889 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.33e-06 SB=8.26e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=0 PANW8=9.114e-15 PANW9=7.812e-14
+ PANW10=9.1326e-14
XMMP0 OUT A VDD! VDD! PFET L=6.2e-08 W=7.2e-07 AD=1.62e-13 AS=2.2608e-13
+ PD=1.17e-06 PS=2.068e-06 NRD=0.369444 NRS=0.190278 M=1 NF=1 CNR_SWITCH=0
+ PCCRIT=0 PAR=1 PTWELL=1 SA=1.842e-06 SB=3.14e-07 SD=0 PANW1=0 PANW2=0 PANW3=0
+ PANW4=0 PANW5=0 PANW6=0 PANW7=4.464e-14 PANW8=9.114e-15 PANW9=3.348e-14
+ PANW10=4.6686e-14
*
.include "NAND4.pex.sp.NAND4.pxi"
*
.ends
*
*
